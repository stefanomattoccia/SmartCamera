`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
X7122ApLy33XagaU4wmSvCY3rmhDYmGsdu52JzcG6DLAV6r9nef79VBnRQmq1ZWqVr/TPBVGWM6T
jHiY/Db6LQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eiWQCREJToriD5/QL6CvZY4Mhm5s/CivoQ2hPT1MRA+pKEJJZ5qwDaJbGtdZNbo0gGIJ6dXaxOgK
IT5TDk6eKeI2RE86mZ8mF4CAM+H06fopV/nxk9BTT03gJLqR9Brp1GS+DdrIR/XUwmjMR+Iv++Ns
MBZJUnnRRdO6UO3Hw5M=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hTGyUtihF9r+b5OhkWCzyWDkdjvOwr5d5s6plhHeCMdFGwzqXyQs+Mkdgb91nD4jSMSSnhqzCiRS
gt825DL8hP6gQRlQmWCgwv7Kz16MAeNQnkipOOuaSMhrHzZgfOlSBcf932f7039Pt1ZDJiSjkJlZ
YzyRZUhV3WXvKtNzxKI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WpFS70W0Y/VrNfYCXWRc2KC6V9s3xozlRNMEeFE/5LLYh0lQVQRqSylvg0/m/Lfzvsxdj5WgMbPa
niFAchkaQOMrbdSjwZAaziTf5IKmrRvz9I7kwdbvZMXepcADpgnDvIkfXzsdz0+tm9nFrjsZOToa
vwwDpESP7RxXxLP+M5d6VjvBzXhxgNDddc2KBEc0QorjgygCd1IMnj1ggE930nAEO9AUus3ajAwc
Ze4wB7B1lljfsDnZduPqvXUFmDi2wA49OPIk2/pa97EPv3pXiLvUtbGYyh9ewLws7hgLLp57WqmG
CnSdjdA8we0Fvt8XF3VV6JZ73LmPYBsY5u6Neg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kYFQQk5eYPep3FSmSvh4UZ7CPdrYerlBOn8iJnrQaukjrQm8OIPk29ZcE4G3t455cPmAbC+JzqCJ
e4SM8tFcF1IYPD/nUGlcg+5TILMA+lyO+v6eiqXLrduWhvgJC9CDW8UgfDv20xScv7n6cL9z/mK/
hVjAH5aNIXl56WR8oY/Mx1Ho+Ojts3csR1iPyuLG5P/eGA6W14BuhOxwcA+E/pr/cJBTTxSIk8nL
+ldyFHLzlm6C6bLKfIIVLiTfag+Bw1swKKmjfMZ6AqHyjcqwWCxXNdPPcHapbj736/wzz/x/l6Cm
U7dDVAkYDFV8g8qMGQ0GKQFN4YU30hPhSZWs5w==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hCamOPW8fbM1ML+ms0Fftqbk/KKcxX/Lj1owftUF6jCvAi0qyhzRo5+OcBSGEM77nXgLbD4GAio3
wV1Cegipn47uDSc1qH2xEFagRWYxXiGJbktPEMOiRVMS0VoIysgmwhvzuV6ZOqwBPXz95+I4sL70
nkp0foBCi3hW/BDZjv/3dbCrmaxD6trkG/JZTjnrgTgXvQmTBwqU1EZ0pHWxMzDRdfjeAj78gTed
JGOAAAfeZZnzLwBdhL5SWhvQ+P2k/yd1ZoMfPy4PM5ZRuYk9v2jLlWTVIv6gj777SWscox6mVt+0
XNzvwTagNjteR1oSAVl+MKwMk2LS5jy4cSRgbQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4960)
`protect data_block
x1JN4qJ5tnTvTxZL3ZB4uIFMnMhDOhHJMfyNrRVvnhzsh7dzZx28sf1IwYuloNXtV+NrbIqpc12A
44gbLJKzcUd+jV92LGjtQ5Ex6TCcyYVyru7neoDhMmSmYAPP22Si/bCJfOGwh8ih+F5f2uHa1kQu
ts/+ZYoxyOGjg2li1NACtNhBvAN1bMx/GjJNFpIJNOyXT9oj6NOvk0N0PAIxd3H+3dOI3JLvy0u/
lv5z8+MS0unObUN0v9LveNrxVDns1LrQVvvMZhI96MFzp0OVasEBTxok0lT7ooay13vJ0FrdwXze
+JW3FIZagk6we5qDsfvAolMtNbHDjJXvHXLpWPZergVLcuhF0oQ0hdXlWSlwbU8Zg5Hjq2iQJXJK
iPiLtPiU+J+QzQz8T8cnT6E+Hrf/mfuiRpf8czIOHT6N5wS4drCBWEYuFpva+Mi0NKTjdJmnJvPJ
KqpwZkuO1xcEMouOe2qBrvjcgBblBVdH5oyfTnvZa/XLTwkLLzH2karNIF/pEHvdb79uA783fvKB
NYtxmtGstdPzkFtP2DqbBA/Ii8o+KjucH8RB37vBbLCxt5C6Dw36yU5HaC/GrgLevtDc05ZC6vCM
2n5UyvzW7cNQHmOzD3tM02Ex26q3siaKN4kfZwnsn3J+tdAqoWN9lIbpxvoFEAjuyNq8T9SslqQQ
qeFiQb23O6SHLH8SuLmEtfUT6+njQH2PLHFysqv7Lai1DOdvVLJQW0AdNtkyQbDSk8dvptiWJWG7
hxNLdPdLfbt5GFF7hED0TfXOpHlVzNxGCfmYYW8La9SzalxN/bEbj83j+f9T2XIu6pDPkAigEOqg
4cQQIh57ZzAuMHibfouDKaPnPQ1R8JXmHTgJALarDezzH2RPysQvljhKHTNjrdHV5apn2Elv1e67
XrPN4F7HlrSD/xUAHyapB6nMFtzxxdmQ/9Vkkfwk3bO5voJ/vdTQKlc8rHE0LA+y6NQZf3BJ4XSE
smO8nNLMqLCC3tuPG8O0A15IifW6txLCcxYhEW1iieAFnM7NVa82F4BIeiYUGXEY0KBfC5oIZHfi
SG2vmGHZN+bKo7HY2SNcMK1645q/SxOimpAPfz/K696shvbcvnuFd9glC/5SWhNcJQCyJyffh1gu
SxbbCMKQDk402zrjm6WWz0MZG0j9IOWKP6/yilQh9cdMa/kUBX2SJuP4/P8CUv6vrJXoNyoClnaK
tD2maashTmzc4/mYEPRLjI/6as6BGw3JLypHFpYlZ7OCxzHVnIgmp2kCnjVL3QdeKffSNQV5K+8y
oJBjMxDkp370bQCBQAmW+PpBcytKEHo4HJJ9xeh/VOKTWltD/IcXjGgfz04m/9NOnwSgnjUGZkmc
i0tMuN/zksAhnExKmjBF2WleSOEp/QhEGuiMlEX/F4pYxiKgv3DEYiC6rbUwSYgjzJkstrur+5N9
8mwrLl8nbCkRGa722scPGpOji7C8YC+6WROxZhMMi5DvqgjzvW9JoCUeX8zAAORJwM4NBMpGvKJI
FGi1LRiaC00LXvCATFq8eGefKTbTMp+TVAg8E64kAwLUMKZ2XTybr10deLCbNhA3YKVMSPukw3XM
L7rXK5RusY5+dmnZJTn+WF6t5H8FmTzQJFwBNv/TPa4olW96DeeglxeoTMH4pWUYX7yaFuRz0bA+
k1FMJiMUGbGo6Krhs1GPMin+kQMyYPKrvJPa509Vdl4kL3+Il4pW/+Mz9h/k4YPXAHpPGbjhLJbS
TKes3uFE929PInrLihczSP6RsWpdgfEK3XgzvjpPP4skoGvZ5rTVIaQZoqnIaIlRTXlsK7uv9fid
ufbUFrHaU9+6Atlt3AFLjKGShqJE7GYsGqAiJTuetPCUHZsE9PJpnOAqjmY3sKIqEIAFxBIcaRU2
m5pQvRRCsDPlDuMWSOGr/apCAv2NBL7+SLxh7HbJ3nuchz01JGT8D40/mRaXxn9bX2mXz2J1MxNE
E9274l3YpzEXRBdyRGPqA8dLvm11JtXAHY1lUwC7pqjzec7I1+krFUR/aWZwtsMyrXTqpEf2FpMf
7ygEcltWEAn4FpjylJIFbIzII2tG4An/sW3endVnfVpm8vma9LTb77d9tnB8L9tB4ikpdPGA75bK
/Jdt3wRgNfWs21QHb25Jpj7biKLBN8CCGT140fWAGZAqyRy9n5UdwG9qsNuTksABxg0uJPV2iQbS
ll/XktaZkadq+3E2v5gEhz4l2tCDiZneXIk7qn2ImsOwz+BdwM23LhG3UZTC3yLCF4/YB+WSyAXG
2Q3307S866nH1nZ5alVzvvjWwzfKf97FUzDBW8vSGJ6kRlk1y6E6jj1W4CymLmiktZjTHpIv3gXb
3lB5lWVMT7OjuOYiK8mtac0HyyKkWyRk+avDwEIXWJamyqZjy3YLXelYdpjmsALwkiVO3KXwUlIG
ie7GXwSfm9HK9a890ffhdDfRh7JLIKB0BL5ImP8wOIovTRHi2lV6/yYLdx05itZYYuUabf7Zjhis
VLlgpCokNx9AIKTihiTqHz382OWaFKQb6ksxzAEMt5DsVFM75fK6hyPA85Fh17hW+CV0PuGifbdi
apkD6BdfVFOxNbd6K/9iF0BOYK+5cuf2B0UuXxiqeLFCR2yxFN099gCagZBtu1feYdqxwA2p+68M
+tW27G06Jy2+KtlNP9Ck0HuYDiIyLSOpWjWDfx6BYpkzmPf2uusDyxQ+g0Xh7RzZUdcx456B/TbJ
nFBraHt00i/UV3Q/F1+oMA5XAHXNAcDEraQe5NnWXbbFsjH8f793TN+GjKx2QaOkr61QTzWQ1NuI
Ycvw4UncZ2zCTfSfkEkWRf+uQetuxWH2tYxNxk/3CiOK/TR3ulYsHLSnDImhjJUK3kWWaRBSBYuH
08xIpxEcfxsv19QVCwnrr3KDzuJxu9LGIX0y/qUnCxDGQxW7sYkTgNYozabxATKTPaEKlpoQeoFa
f2KSTR1Q1uetMO5CkvYCf0wVa8uhhllw2TFX79GHerNrmJLDDDThsRUF9wjJ4gEUiawAmFGE5WIc
WEMLS6Oc/Pc4k1KYy2bIQGlpcdfltfxdief5olEA8Bj79/ytsvmOSaXct2epoaYYS6FJUMxT/ssm
+EOZ//PbWjEb0UtrauLAqnxtDsMSLz/f3bJx+ud/OI9wwMUyNVqC5fa71nPZgbrO8xtvOQxxbuyt
uVnegt8Wg3dG1zp0FTwluNeKaqKTDw67c7qVhLmlKPjGyBOQgEUwMdoWJn81REnjkk+NHs8QvmKb
1yeKoLZMkEp7rsWp5eoEjFU2ko3uAodc8D7OCaR6JUpmZ22N+/cL0HkbMU2N7GRDBBCrfLq5zO13
ZqzWdkxI2MZ3CdzSPSrxems5WgzS3iduqlbHW6JCqA3G+dftxnrr/2sY38Gg6vVLVJNenSl84KpH
Q3fLoyKlcGxbwayPA9JOPZ2MfCcZsO0VcBt4o/LMSMEJcDFZCS09i0BZ61HOI/Sscs+55fvyd7iR
GYofVdYOEwlg1EcjFf7xinnS2L0zGoana3mXhDk5oe/mzuuDm7850d7krqrZKMzSWvvCTZvtMXZg
OhhSc5DGWpgyyMlwW3knPO35bCNpUQo5r0Rl61o3V3aldBbRf7VvASN+vw3WdX2cWzGda0sNL/vW
AmR4vgse4j8P2jdNUSAR9UaF1/niEysFuWdRcevg2SXY8fGM3o2tF0G1KA63kSS8Tn7+euVTld1l
3rZogyhUuy7bHMf6SeBOpe8LouroUR890HUxP7c42BcJAO7IaXwEzd2kLF22xsb2dIqrEh/erv4Y
TR1wzQQq03Xig0uvA4KLngwwG+jUIamH473KjDrVz2vlvCX3mFTqOih8Cn6YqxLixyY2VJ2G0/8q
EkuUJIl9Da41dPa5jzZLlHqM7Ex/YqkNiQ827VfyNy1o+5miIT4C609bldfXbeLWJnHFEC6/PF43
AU1nfGCgzS2onN+sc9HEAnrvvBVUd3gIbOB4YJu3JtbW0W+7IWGgenZ8bnejWe2oTogw94efGtpj
RPIufzXh1z1VoJ166HzalxV6OuCeCBy8nDFy9kuQS/6XKrQsl1GCd02Y7C6K+Xc/ypxaH7hsTaFJ
saFx3yKsrHJ2cv4Idjpoj1OO7NmHwppvoGcv4kJ2m0Tl0XjKsuJYzzhSPyQKLG6P1teWAuoqhpgt
BvX7ttY+LsSDerqiEyLdz/sgB6JOgTHrBcly6258uA5hthADIUc5xoeRiYOIbeo1NrM76cn8YGXV
Sv2hDukYFuFEUJaaB7lrxPnHC8BoaWxVbPuwFskJookAScP6D5A96UYTNTIwsVfrCIb9j8Yrz88T
0ScvoBwrhym6hSsN70FSLJugHb1RcR9OFUrSG14GXIwczIxlC30boGuzDbXM1ZnwR5nmKjTHBdUj
EBfdRMsnM7eMExvTv2fuA9s/wr52dd0/CGAp0r6EyApcawKh1bQcfOSUBwiadb2Sa7dabo4oHCfB
XnCE/n11EfGBy+RDtk8xeQDGGT3h1pNA+WePZMTO8x5vrt7UbCIakoqnx+5zNKBNL9O7IrMIGGww
P4yDBIjH9khuROIftmMDoH3TiWfLkm+RMP7H/KnM4Cqws0QOc+ZlEBNnT4S2Q2NnNqrhMDExbfuK
0ZrEoAlMwZz1VbUshl7qYAJNahEFGgfphcb7Ci5FI2OjBB84ymBXR1ZFLxKRU+h7IVj14axEHvlV
nFJ5LENqntmq5kBw1XYdKs9hobg7/18ImKKP1jyMHYyUAnYv1n0xVi/kASFOwol0+il7P/yVpYBn
ehfySXcd5QGDcIMC3e9oLkMxdeN/4Mc+omWKwHEbRZT4o9vcGG1uEn5m8Nhx3QTK3xO59NgmeM7J
2YdUwDKFfeA1LEJ012KxkI0s7Tho9EjG0BBP11mNoIQhHfMfFzwySL2ASCEDn8UqPsyuvchxHauC
VHyXP6fX1zdpd4xLhjO041DsjHBWANhg5PQXDZwCf239TwzmU6GCLTDhtAVbsDEQ0Yj997ltF+iY
JQbywglnCbL9r+ICtEfPVN6wgn1q74950oP/TNF1ItjvR9SANqhATiZ2dhQWp3PeNuffdnNAzk9h
iSeCbhwPPKSky3egN4TFTvgPkhkKcDod5NGOFEw6PIuTW2FuI3EqcAA/+o/JmBh00gK6Dq62/0du
SrbIzIDtxse1OXJ8UKFw53biXlHX6rrPlfmTLHjEK5eFw4m5SLVZR+SLt4rAMJZx/xrgISkBXST5
AA2mPG+gW36JjRVXMYBCAxvg0J013z2elew1fVdWoz9BiZEF3wfAHezxg/4bXsIjQOyb3W3n+Puq
0NiOXvE6meef0hOCjGhKHeo/jI+D77r0yrbiUXm4R87yRxCBrfNzjMmn8JtGC+FfNnT0pFKVU3yk
y3XMQJO23kF1SgR7DD7X0adJ/KxD5XLP5tB06XkXra0x/l13+HCTEr2eaQMJFnYcGVQr0NW4maDB
iFYEGqHAFohham04EAHwBswQK50eRW1CUtPYfgZ83Crho+12Hs2AWRDVIzyYyadnze1UEM1Mdu4q
NMWyXuJPe7iSRQX+jHqJBnYZnDJjqukjfhqvSAAMY85T4F0rR8y4zeIail9E8Z3EiOSF/F/NhZ7m
CTg0v65KY4YCK1omwoklKWUIqvp7XIk7JFrCGn1FjKeoYvhfp7ZCEF7bnMQB0Hiy45DBF/hfbFSp
0TgIn397lSPuqk9oP96GlMwVh02YpInZass/Baz1Px++tFhSPBJYXBdemaO+W097/hGrVaxCF5+2
7WjR+wiLVhBx/xrIWUfPnw3iFoiT/wu4NhGhrDJfCG0vnnNw+9h/zFnGisNZ2+DSE8H6GdrdUowO
rwNGEqDBaV8QSdjbRiCJEHpAExB7sWMkSNCVjE81rF5qqoIy+FYbiZ6g2CXskRJ8k0TEAjTPcp3e
fx+gH+kItNcPynLUthyOGIMKq6P8n9kQCG2HeZRaAu0sk2ZLyILPv0qmODrpDQPDjvF9UBKkY3YA
aJHusEMV9xI/arB81GJrxqD2ryOX7C2iIcbFgiIIyt0tkECE50/Ui1e5MGG6/4Q0aQlyexmiiDy5
AK4g0QVhopCmSrRJH+jZ/ENmVBKAsNvJTv0dcfogJ9JXILHbIIZqIAeDtgmQy1h+zQMGlGZTGCwP
9czjwxlPEun2gV4VZBEmhb9npkDjZoVU6ryh0J9uIAl9avpwo1IV1Y6+/izlipwIpCGuXEoGESP0
xiY/+SORF31osAmOUaO8DULm/+KrEbX98w0GaMU4govC6yTq3nMgr7LmNd6v3i3H50RxUerowwJg
fIhGzSkfVGYFQagcSk2/0UK5zGpxCyw3rltbd34ESAhwB/V2TyUbwbUzkvrgnTv4cunOaZCYyUSQ
a41GOkxX6IQfn6OPaC3/MLDWX4BUU0b5loBGTsFNVZA4yGsyJtr9cpPh2Fe3Sxi97QJH39XiLWI3
LCvUUSJsMLyiONMKRdIEeX61XUSKXG+AaDZqfMCYwAI91kM28Uhk5E9tSkm2xNa6CFqG95NLjmUR
Qw5UvpmtO37QG076FwOfciVXvmilfDd7BACJ9SlGdlrHpdmkrtBw3F7JFjGItFCVS7hMiK7pvg8d
dg==
`protect end_protected
