`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FEMO5gEygrepbyTIAb6bnTzXzKtTa7hkErwuF8UlttB0u+dyJHGgNZ7crkojw8pXdXDcfF1p7dA+
pQaP5/BGSQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BUAwVhxzmgAogQkTbbeTYgQQyI5Ea0fpFwP7NYo/fJYalzsEKCNo+mHLYdEEN5P2wAyI2jwL1Ldl
2cWWTvWw0FFDx6CAqyMZZ6MjBcXKMrbvZz5x1XnEF9Yq73tmyh83lBHL1QeXvwFWsV/MtPawWibr
DqrVdukNDMYsS1phrww=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S/0xh+8q5ei48mqpxhA9UHAZBmce/qaAZdB8DypuX8HuxWaop+hJCz7/amofM8Y/1RIn9ynwmPIG
lcSFISHwXxQw0TOGzhwmVeIUphOOW6Xj8efDxrEsgqjlN4uFDONpJWsykX0bjYlxDKh7V8VYmxsZ
W2QII8Eg9roJuKe/q5c=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m4EIihJzHXIjlJlX/nPXOZoP0R5PF62b4QI6DPL+tjjKUW02RGUxgKdMgmE9mHps5NWzgwv1KD8/
U89gIWVIYKuI7AkCRzSIq4+7kF2eDJ/Rkcrj2wW4xn9mJfkpoCsS7AtOGt49NAv4zZwBC027t3wc
ufboERWDi1EvdAKPgGQm9PlsQcCafLmx2ptvdo46UvpFqzYZ1W6ZCuZOinFXuDbR5Dl2XITXUKEf
6Qit/856vn+C1AiQMPBPg5t84jX1T0muMNdiJagE6NH9TuIZh34Zh8xMpiJVMleWEJ5+ar5ZYsLd
r0bHpLmOwwOHnlbs80+gfl7gGs5ckUJar8uTrw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ugm/yKAo2KdQRz7pCWPXE6yTuk91zWS8vqvbp4N0Y0rRLeVjfYgYNsoxanpin9oKBWGqB/EwwFiI
OecyJhZzQraiaozD95T8G3Czi/CyjQfIuIxyZlOURLuKQG7CmONNSV0/exWSPuBfn3Pm6VM3OjmU
JLfuRDs2d4YDFd+q56oiiHQQ8vCWNnabDnJXcPKxlSBuxC2iBafhs1u9xdnlfbPeZ3KQYthd7ZgT
hC+BU1U9gXilj5HY81LPuP3oaZbJJceer+0o1dASuDQYfcDQjic35pfjZvrWfHg/SGJYnP9rBSDj
+CEsTamUhMcogvVE3I0C8I+NXEkM9BpD6lpS8g==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QZqM4wdZAFPtQs4YrlRwMrWNZIys0rSI0ZT1kN94aimnqT96e7hJXmu8OIn/cJHN+QLJpyX2bZsb
9aS/bO2EpwxEH9ivoPATAnDH84ywTGBY0z4TDTpMdmLig2F5x41qoVx7Xjt+NiM1WzZMdOXtb6+T
7rMRng3bWtMuYeGIO49nyrXfIsdW/BWSAUnc7REbccqnnz50wxmKOz8/Cxc0CzxowbVvovJtn85V
3ZbWUq3enzYLdYiG1rbSQDaPniVAqH2+PhUK2ZHB0HY/TJkgvwTPZwQdfAanCA/ekvY9LLeNdJeh
Tfdqj+WcsCML1NkALEeSJjr2A1ERcuQwgDCfyQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6000)
`protect data_block
VfzJhJrgqQcpoMLB9xda1JsG8+jZR5TLvYhH3JlEnCbbeGJkX8vN8YhLaPsfk048aKzQWZqzH2j1
JbY/bUAEOtVqxXp7jgYhL9S/fhF8IQorV8O9dILW/0mNxI5z8dRtQV69CphvdHKJ5uDipt9O5WQ6
YPyLCyrZigPnRoRJrgEVy1ZavxIj2MZXJHnfFxWGC+80DIS63pIi1jvFolqGTqayk0NB8CCye2tK
7Uh7myhZzNnYs4d7rmF0SMcniXBQUxq3OlpLO/KPMkbD0tGS2coN7TmKbqmytHnz6/SOTjSg2JKD
/iMLxPO31HuN+x0v5+/KxC2O4KehDcWb1LEfb6uRAahhH7Aheg8XICA35A4mmDUux/N/uCPQc9ZB
VwdxdxmypQnNTg3aoYcoVqZvqst3tBztVH04HOEj7RfOjNh2I9hveLwzFG8hXqy4sQhFjD+PSNzc
DDz9zAzbHQ5GjuHf/reEkEFGLzT0HG1tINvzwE6Z0n7biBKnFaW5gmzjqunmxIVAWglIimn90bpc
ZtdHLiXRz1ejud32UolaZ8FPO2M+Oh+G4LZKjpu4Ovs8M0h0QLYKDvjqW3oiIo8FyGTK2LMeDd3q
W6qINUyFpvHvM+F0vGgFPYUqL/Cr9yl+mjw8LYRZxwx3dPYe9GdNMixM29MyobcoNYX6LlnZ3lOC
QLC7yE7hX/2EiGLY04z3KE/SgSTcpMDqx8dCKimwi6Y0JXt1Bp6pWs9UnKK5Zwx7/M5cGJJmdmUA
RxUmQWvRxLjsoqMMW34feddpqHipmWfpGEwwVuXepvevWR4H7BkT530kiehoocHIs396bWvKEE+s
BK2xDRH2IYcqmzBH//ZKiwFl82h8taWsHhwz18o/UOxS0D65uKav2p4zNRbl+DwXbIERtl28TfSu
lxWXsZPYyM7QGuQDRaVTkhuf7vZzcltUkvmPbIZPl4mqVFgCQtKT/qrfaeSm8gtm80WXeeIwSmTT
Iy7W72vWVWMZOqYv6K3OnpHR0xedradyLddlJ/XpBdiMJ9QM+RlkusXjIGSAhWfdpqiy4GgNFjZl
Y4oH2ODfE6iVTEwO9LQu6Zackim0AtuaaTdQADshtFFF3ICZ7IOMqlFQiXOdgW7cbNFqb2JR15tK
4RFYeb3NYRehUL+TPLx133luAuM18r1AOerI2sz54heyjnNjMj92LemW3Fq0SrNa+9ErbsWZO7SR
+0VSqXjRSHPtOGgtcy1PgN6wszyMchluZFBUHvi0g8D5Fql+kz7avBHuS0z3/qUfBZ5WGhunuaPF
4cTcZGN+aBvLSIQQskio1g2j/tdQKmpD6e+++yLL3IoDp/QqL15F/b3SXg/S2kyq5wfghHI3d1lx
42REd1D1jpoe2jClOeIRvpExNunBtq2SMMF149qXurDoUPD0TwTHYxTOdM33cz7g8jWic3kRTjbZ
rN0WfS0vdoB41GnsObexp5WxH7F4tvzFG6eCLX3wfAmsU+tRpJNj4s/PKqxJimmhJ+DegjToyTjB
CSRrCz8oh6EiV/XIgPJrRsvIvfFAwBo2kX7/2VKa5Z+ihRMs760let8ytSNa5kkoQfSocsRMjfLY
PnrzlyOz7+nCPCAEs1OhKmPkNIHDFz4Xo8GRxePFjtIHVWOYY5F77XyYWnQwV24Adl8eYz1+zlkx
am3A/Am6f0L1dWH4oKaBVfxrGhvfsCXZ/GTGSfvw41Zo1M07T7XY+Ie3AZacTuW30FiKqgQ0qDmp
pvfTgSyVAi4ZRRRtIMXIB058AbPD0gO+XcpwzpJKplTZ3gLo/8KpGeVYrb+41SwH3Mkm2NORCWqs
qOjSufojqK2bN+JL/6rVfVC9SvaAjSjARzl2ktfneFjH8mKQAu0ITyP7pxXy2K91LpVp5i5EvAHR
kjQ3zBiBqDTmhVEyYYOBar2H05OuT2HAXdIex5rUXkSVv41P7JLLNEGB7HcH8y68SMEx+yEltIn7
PWQvu4xE0EWyG44WeGi9EFjwdx0LeTYj5HPGPiz014EuJL8+yIGQXLEpRQTs+YhZ8+rdKBUvbglz
3IocuWRdqCK3WfXgVHvZ0PM7/HAJdfvYRLi1MJz2HPwG73nso3d57Zg2BA1/fqrjKWxFkJnwpdEt
dn5w3mwmLrlnEWod3/l/IiRdBGoR/fT9Kl71ZEAtQ9zHT2wSonpsaO8gBWbNihzC5ZDcrH5N1OLL
gxPYYICjirKKUnTelhVR8ZITWF2yN+1bRj+pCq36LoagGRQIoo7YSfDACmHL6Bb9jVYU46Ki8cXV
V6F0R5hL0Q+0Y89XJ+RIBJSUmFclEd8zDqfpzvTLgcGETG1wXeY8NfPZ1l+JEPOWDlD3kwDzREil
PUtD8unLypE2v24+aMMV3HJbsFfyh7cTj+gIxbj3Jl8LuAKQ7+ZxulTcW6mIg8nIb/9i6JFuPWkG
JVjYB7WyHpxkr++tRN4XDpSPlydO2kYgqJs5swV3ku/DHebRS6gTj4UKq6H+32DbQ0pdAhIXfUGa
95XzwU7Km+VIyuEuUQhk9M4envc01SQt9nmpAaurM37WK8WnwEYSvhLgsiwniKoYE5kWtPCNHFiV
ZLkiOlPZLApXLxrDqfu1krulshGs7YocxO43ABSsCuz+g3Z3YzCT26hQt1GB+7xXwpQblkKgBfJx
okyzKeJA/NI3pnPDLMQurpGn0+W6zqVaJ4X2JyvSRJSjXYtylyBz336fo1MYVtGNg+FG7jb38iPg
Ln68ZHu7fKMPptEo8Z8mUNLxg/zc6byEnz0TYF2lTrFxexS+IgoUK/TEUWQCUQFasxwUzvowjJOi
qlixhV7YBBb8hdKYyjnAG/dx6Ku2Zj4WVVxm0W/giID2wrSZ0MS/s5jLuTlGkaHW0oWWddsWKm7w
2dUUEejtD4YCD4kp6NsSL9+IY/DHSXS4FFs04L5U0pL2c6h+ocF2ewvPuSoQjQtRfUeuT0gN4UcH
rTu7zkkEp0PwLKcjdzwKn77g2kwKSQh7i7WaQ7wILDUa7sK4PN8EVgBbT79l/v7nbhcKQgZ0RZiw
tCNVN2/nkrLAsDneDd+O8OBFLFTu3mPBIJWDfBhGqMpzK/DESS8Cq6jF86AjLLUsNOvuKVXVJfo7
0xJag1BRRw7+geuk5qQ6QGsVc9k0V5UzwwgfsZL5oVYP/RMoQV5HIYRUhvXqdfdfYFeP6aKi3He6
51uMLMBIATrdG0D4aUh5vPMkH6RKsguwIwdg19LhilZO/jky8iziukdiHgD8/rV4hL5Huu7RW/6r
B8rjdBiGZXXwpuDPsjd1ak+3Ro1Ndw6QRBV2WTmXwND7yMYOOZzen7BTihqjg4wvEvdTiRn3npZ9
VEZSvdkc9hEW9i9dh/IicwSEDZFlrNaSJROCuRUbLLHWlhz1jx4QuzcopX7542m8ZH00TqB+YtQn
LbqbpDJxXGj15j6c+8LEqgmB0fNTZ+QuEzHidx7OWuOHWMPsA/gyaKR/B9W6tQpnCX8XmtcOIhEF
yaXi5gMGwxhBt/9vrBfA52ja7hbQMd9iMU89ThPJNLz5+Dt2ukWwHHqFt4fGkLeHlmyHK6ZH647D
NWlIlaaw99jRThtZnzJf9X7NQrq/i3fE1Gc6osvOQnYOhxt91EAKjg7LBQquXE8zkoGDBijJHShy
SJwcuFvt5YR4KqJqiJqPr9CJcHJj2oSl01sjVtRxaEw8qO0Pw5VWAqDWf1a0rMuTzltOwlJmuUe4
TNN/VdXtnxTnIHN2fr+BE7e/04d/gf+13tQssU/mMW3lQLH2gzGdowp/5mWlju+mYMc9Kz8CcLNp
jNJVhTSocQJ5Uvd/eZwyX/+aPHw7d+lYE5Ru0Zt+ciyIRK8GamR0B9CfDNsTdIqGeTGQRYGSJTog
FcyD1lcZw7VAPptaccPajvcsYJSU5FakfQ9ONyt6aN8oHoZTzVUjHe62zXD2sG9Vozq/CV2CNWaO
RS4syE8VZHJr5RAbxhgvWF0aCZHko/oLjw4LxcDonyg9+kb2blcwDk8BQnRQVXrGgCTCzbRLXOtU
WaQDMlzRFefA3MsJnTcQvG0PH+q+EylBtCL24V3yYerV3bvACNXYaFubZlpyE6X8DXl/uZ3gHQNt
lnE2OL1lggb6nttyN1WK+2tk4ppdc0yiGIpR5v4wFp1tAFV04X0QsEvHwK9RQnbk6LXWfpQ2G3nK
gVkZIG03YqJ2vZqxb46ijPTVbbdsI52AjrQnRbNt8DygfTSDrarK+/My892CkyDZZCZVfsBoeanf
G9fiR/4Nj3xZMNE2NjWuKZKv9cmqE9DQcAOu/54K99Nha6k8Rh2KAJzCmgX2VZn1SFn0CXFkV2ef
OfLkP4ONChE/i/xcI+72twS6PsM2ZtT4gK/vjZfRN2HojhkmDdfLeETD2bq08JeGzyHlWorrcZA6
+dEP7IFCt0WkPFldJ2G2iILaqIKKAy+sUBwa3fmfAvOcixxZoxgxs7SjcDn7sRShQhGa5iZ6ZVx6
UJ9Yc+D0eBvs9/kPrAbmQJbsZiS8WfAuzg+bt6imcMUXYXw/PLQeZD4TJ+O06zlyCfhSvWo7rVD4
30E8HMO26vzv8kbdvSwvhHfvam8v+Op7FxYxsbSgWwURl00Lr5/9EeadDNLaq55NIoN2fb20pBs0
QBBtDVAxOxTSp+j8f1+DL4rzJ+7b4StponMs8u9OnDJiiX3vzpB1TTXbj35G4kW5fUIgAfD33byD
kGI/b2cme9u9TW9VKjgkV/obGmkojd/rWK+Sfb9g5BRqiAR/0+SrYDemqkn2MKPBCaHp5DQ39MPs
S7rp/BMeHxxVQjzOsyrrI6y543EbqM/M0qjjYkqATw2zGpK41gv7WSsz1byBm3BuBsw1onyEYlih
9mhkzmOeJmecG7SynF09fcU12Yvzk89XXSnMGVbmTPaSr9ryxjZJOq0rBg+YrC0lH2MaAHElPxxS
NUcg5ThdQhWjyGOF5ifjx2JJHILZZ4+4Mw2RsIKTp+WqH1srLL8BwM4T4219U9tUnv1r5dkPbn1a
bRpF+y0buSwOsjibotLkI4rAIskoef9NNx8SmAY0De8xCKAmHAJooaneE3mziz4i7jcLH/UAmoXS
4qJiqOLsLocw1L+XfFjBuntWqn4xRIkMSN32CkKRfFlFBTrlBfm2vluhFYfs+Nt2zVFL4w6mqnS4
UuIfV+3QwcDiOZfDfc/qqPwfdnf50nZBkK+1+baEYAjolrhjdLaAHKZLWmoYRY4PDTTQobcwlnYy
sDGBYrtVuW6NR4Qa39wiHri2MK2Dd7pd5EQkdNoLnNQIf8y8GW+ATVYy56T5JUGJlo+CCRymhsQS
b4JmqVm28B90GUSdwyuMqsWQ/63jmUiMhEsG5wL/A3Ux2o90fJY4ggMDS0b7Jf0lgTAgpedpJwvH
uUVEkCkk0A6862bTTI16KzpbAyvJMEMSDYDNZ9n0eeFqLORgHoG24oZdbhE40ZO8LJueaQB0nATc
cJJRRlyHm6a301qCjRbquW47Vfi4CgOetOJ7oYfHmjjKPr0knsajgrFFGIygNjX4R5JbcsRlK0DG
JlOTvSQ3dtdkMg6s6ilifwzxq1nAHnEN8pPV29F4frgcS9EK7hfahZO0EUYE66AKHsp2GBdLYLJo
ItaUySNn0rLXUSegEcAKsOTDDtcitzc8lhfONs/QUg0SAy4cXehgghU9D0DscbUwUTF2iZY3AHMz
4MHGB0vP77CuHEC8E+z3M6SYabHhenNRrQCEFKkOB+yhNRR9+06LvcbucqsgUsnTLXQVcAQ4iD8z
E3yfecatnrLiHc3p4Aqh3z/qoadWn2KY1i2excpNZNZTS8SsSirPRrrK1vvEj2nCOQrOoSfsIeG1
hvMm5veJOalKpQAPVpkJ0BuaWbQdpJz/LhTfcyinC7PB2HrdFgT4aDz8DzngMUhjeTMDGpNIadCA
xMMqG4aAKMPGglgu80C4yDauGfjN7NFYvtCp6GTOR3Sqkc/0BvWKiyZhPrmj11uoM3uu5CHX6P8l
aSNsjJHiUgfBs1PLDe8D9Otr/iJxzc60EPkgDOb4HTBVO4wABexw/t7g0zVz0LaVJRJUdjo5fTd/
h6ZbbBnQmRurYXlQfj89cZr+4ZXwUVvr0+ZjmN1hrxgraUWvrPC0WQvZLDkZIjLmJrL9TtJRW9M8
a4GF+ne4r1tJlZ79xqzrbFFQXsRFCOLrcNornNUO6IBeTGCJ/9TSBKaiBFM9cqL1KbZPOJxWRRsT
S+rGLpJuRDDxG6moC9ZSS9FbxPYVatXXsrosy30eSOqtd5TOpwtWigs7JdFlHT9r5W8upCs4yAZy
IXHafxlV91CNt8efufv0IR3RZhZxLULVUKAY0VZ2YfOLgjkrjzE4ljU2r8hXVLNNT8As5M3Fgstv
7YZ8x9uHaeBDCYLejffJEPR2ArNQSas4biuJTikZEFQ0fghvrEs4SerzZ5Ve2n7taWvvso2gEVVJ
SFptuE/KfoT+wryQEe8TnmE00Jh2JNYgif8xASPlF3UVsGzcvEMrBelPhqZlnbZAaMxcT/PFMI+o
gwTKueIytMZ9q6dSB2+Gqa6+uHj4O76nyqrLTx4ESO25KtTvI4EcHgKOTtDPYui16m2OzWCSVzG5
8R3zkS/prrD1Hs6G9Ejkmvel5KmZMM97GUuqcHdw7ESDemjbGctb/YV+dr7F8ZMFFTaeQdddw5X4
shdLluQB/dXBcti8TeEv3AlYwVLT6pYoh5EFlCGbci3wwpoBdV+4FZaJIDLyvxAl43jhMtR13Iqe
dS3CKaf5DnSXftCoppYV9Jey6fo9/ufFaPA9cXRW/sExYppif/8RRox+o5FZNQcyzGfpDq25AU2/
nO81OJ0+HMZEk5VnSxbh/drwhCsrX/9Ut0A4wu0TAdah3JO9XV6u1T+r4/wN1fAmAK/NM//F/tRz
hdLSUn6oTxGQUkhMLwMEoYEdiOHPsKRfi8Kxkr42Jb1/64EJHbwP0aRcEzIeT0NiFTsBiQ3eurtd
6yDVjV8vxvF5ZXtHTUB7FNep2Xcx4SnZ1Z6cNPI9/apFyDb2tMYjm7tX+uA+5JLZnSl448KznR97
6lSOaYNQADRKCT+pJfSOhD30OwERD2wulB2So2ljXx119h5qhngj0hwX27Y8PSMh9XJDEuE2qnrv
mzDcM6xZEKOsJ72WubsjRPdx6d41ZxtDdjFsBZM8Ig1zgByhv/W/hc69Isr/LLC45XfmV9BrXt1n
RsWfJkeJT1ij7w7IaV787iQmG2eoZ2/Z070M5XWSxH58WFBfmnuZAXvogN+Ku9eAGWtW9mklXo9G
iKbljwLq4hVczx7hAMDIxKs/6/CKTHcyJsZFvyUV3Nwi6FO8tUYiyDvmYeHVtrhjSuj26wmL56vA
RqntOP54a7hvs+JUzcwtB45muX3smWtEWqSwPKPjKv37XRHWnMJa/YK5r1nObeAfKLl9liSuGb+r
0m/KhhNAy3soRiOU33yepoyh4/zKfEl3KDnGYc2uQL20gFvNU5CVxuTHvP22Db+ldU5wtnEAq1BG
xHBg9YNU3stUY4q/SYudNdoMvLt9KY4H1lmoFq2IpcIVTU67U20b9DrMqfvBf5GRZUcrp55h8rPK
Teyk2PJEox9byZDhoDARWEHrvSg0V4xaBDD5K7JYK94ttrwor/5HxYBR9sZUlzYt/ukG5E7kAJSC
8erMUwJIXbAQkRgRZ3+QVqeSpbYtT/JOn1cMz/TDbCi8J7y2tWMmrjszds28posT4q9tSg5lIJxx
QT9hJB1Kd6lPPZFwKK2dLqd1Pr632nu7Th0kO7gyeB8H3TsfQ6Yoi6fFPBMD8cvIFFOoER19iNVH
fp7b7U56XTPqgu9FdM/goTt4DRk0L/eIeUsTNhw7w7AnWGEVnaj3QN2bRrk0r3EpdWDcMLcsSIQd
A1kmwH4aeItcwcUStCoANWN43QKj1EboAa83SQ49pnXyZAB5MJishnDBOhFmO0N17tb/Q3k3Jp91
/HrbtVjHVrlmicUBKq3X
`protect end_protected
