`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
X7122ApLy33XagaU4wmSvCY3rmhDYmGsdu52JzcG6DLAV6r9nef79VBnRQmq1ZWqVr/TPBVGWM6T
jHiY/Db6LQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eiWQCREJToriD5/QL6CvZY4Mhm5s/CivoQ2hPT1MRA+pKEJJZ5qwDaJbGtdZNbo0gGIJ6dXaxOgK
IT5TDk6eKeI2RE86mZ8mF4CAM+H06fopV/nxk9BTT03gJLqR9Brp1GS+DdrIR/XUwmjMR+Iv++Ns
MBZJUnnRRdO6UO3Hw5M=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hTGyUtihF9r+b5OhkWCzyWDkdjvOwr5d5s6plhHeCMdFGwzqXyQs+Mkdgb91nD4jSMSSnhqzCiRS
gt825DL8hP6gQRlQmWCgwv7Kz16MAeNQnkipOOuaSMhrHzZgfOlSBcf932f7039Pt1ZDJiSjkJlZ
YzyRZUhV3WXvKtNzxKI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WpFS70W0Y/VrNfYCXWRc2KC6V9s3xozlRNMEeFE/5LLYh0lQVQRqSylvg0/m/Lfzvsxdj5WgMbPa
niFAchkaQOMrbdSjwZAaziTf5IKmrRvz9I7kwdbvZMXepcADpgnDvIkfXzsdz0+tm9nFrjsZOToa
vwwDpESP7RxXxLP+M5d6VjvBzXhxgNDddc2KBEc0QorjgygCd1IMnj1ggE930nAEO9AUus3ajAwc
Ze4wB7B1lljfsDnZduPqvXUFmDi2wA49OPIk2/pa97EPv3pXiLvUtbGYyh9ewLws7hgLLp57WqmG
CnSdjdA8we0Fvt8XF3VV6JZ73LmPYBsY5u6Neg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kYFQQk5eYPep3FSmSvh4UZ7CPdrYerlBOn8iJnrQaukjrQm8OIPk29ZcE4G3t455cPmAbC+JzqCJ
e4SM8tFcF1IYPD/nUGlcg+5TILMA+lyO+v6eiqXLrduWhvgJC9CDW8UgfDv20xScv7n6cL9z/mK/
hVjAH5aNIXl56WR8oY/Mx1Ho+Ojts3csR1iPyuLG5P/eGA6W14BuhOxwcA+E/pr/cJBTTxSIk8nL
+ldyFHLzlm6C6bLKfIIVLiTfag+Bw1swKKmjfMZ6AqHyjcqwWCxXNdPPcHapbj736/wzz/x/l6Cm
U7dDVAkYDFV8g8qMGQ0GKQFN4YU30hPhSZWs5w==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hCamOPW8fbM1ML+ms0Fftqbk/KKcxX/Lj1owftUF6jCvAi0qyhzRo5+OcBSGEM77nXgLbD4GAio3
wV1Cegipn47uDSc1qH2xEFagRWYxXiGJbktPEMOiRVMS0VoIysgmwhvzuV6ZOqwBPXz95+I4sL70
nkp0foBCi3hW/BDZjv/3dbCrmaxD6trkG/JZTjnrgTgXvQmTBwqU1EZ0pHWxMzDRdfjeAj78gTed
JGOAAAfeZZnzLwBdhL5SWhvQ+P2k/yd1ZoMfPy4PM5ZRuYk9v2jLlWTVIv6gj777SWscox6mVt+0
XNzvwTagNjteR1oSAVl+MKwMk2LS5jy4cSRgbQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18016)
`protect data_block
x1JN4qJ5tnTvTxZL3ZB4uFImFhJ4FfbrWsjkgJBiGnGJ44qAQSARu/5TNSegFyTj2jx7rz4S/5KP
EgCfhZVswjx7SnEMju6DZmAn5uvfMkS8lZlXiGWMJmxGz/ogSDuO1tKDcsLBxSjOia5wSv+KRWsF
t+Zybzp4+QJFl5t69IMS1x/PqlgPzTWs5s4Ggh0xrH3fiibzDpqybIIBvIOocp9B+4o0a/sVr8vW
o4CiABZ0D4S3F1QmSbmFfWbJ4kIwnnjRMWRorQNgYCUbPFSLpfKYeJe2Imm+7qMH/2lCh0t4ioqW
P9EUn5rYnkZGlqHdurmB4R011Jc823W7XbSbesa+dlz56HTZxh07taDpUp9f3zNOZYkzRQWsOAEE
78BKAPyt9szYkTFUbtRvi51wYZdWMmMDBV2p4Ho/BYSo/YatPKc6chYAvqOYRsBBBT9INF0aYiQO
snRmGDCfx6bU373gyka7pPZg+vCrdffCVpVYDFDfOEQniAyNxyYQKAz1+6/mF1PxHocZe/fXa89w
+sbHfiAVOh0z/c/AgIRl4kKvZq1LraV9FBinmnsdf1pqpMaU0XdB1zHXI9w66XDihhVL/uK5IHLO
3IyUkBktfG2rNeYAiko1kf5A3x7cWZai5rWT2o7qlvJmb2iX+9uaV4uIsDVhcLsyAn9gDXb7uWp2
aEhw2FdV/0Zqaoe5/pFUaRmxO3pRbPTrj4P4f1ATMuZcdsIQVTsAb08Tx1/UabuUeau7td/XKFIs
9gj/sVtcQWSWtWHXOKlYZQM4QBjSnZTrD19x3xWmd9ki1e8fOntHn6CumQYZWHlb/mdmLpgshls/
PNNmT06Q0A/c1yvYjxOCVF0ea3O2Itfcl1BIgeLFuu46ammmZgqR4bS8/8JUu95VeHVvXuo3mPG4
6ln86zykXMXF3gKgDuuZDSPyhee+OeEtJmNiQlPgYCX0xEcbumfcUVtGP7Z489nO96SZaW5onGRK
gE5MMkcon8ubZX3bGxyjzMzRv5VD1jfe6lI0MyYeYA2+9OWdbGjV5GCbpypl6QxFYdXEUMpfVFTL
EWBnRPAMqNXdL2g+/VAmjt+nKDOZcfZe/Gez7gKm+9Coe1NqRmIAZbb0yg2cxeRogMyuZbcMOCY6
9wtm9yqyqc6NH9yO6Wc2lDN7qohvsRzJGE7uA/B2Ugdqmkeqzt6DMrGAgYBC/3kn2MKqr7fAdPiE
y9b5tkJxdkxyQLklrYJCcOmfNiqdisfB07aDi5vGAytoYIbPV69pX1oxtLwcHSdaoNDTJ5c4NGZ3
kROzzmhfe0J/wkOj3Z2SdOp1sHehBIkOBDkZ7WJ6rWcBFAXZm33UWJPjclQXPKEHZ5wpQm52GVFl
HiF5y3RW0Rv9x9rkMaz7IJVrVGv9W8KiBl2IyROZI+LwLUPSMfUAlcMlAFLcNVT3Q6b6PcDpaLCG
EhnuzHUPAZst+mdiIgCgyWz9muqcdRH+DIdCoHGSiYtEQ6hDrQ4NT7SpCZnTyWigR26kOoO7SMPd
p7EMAE55CQEXr8kNP3xM6WUlg+ov4p/n/Wp3u5Dasz2OdkZ/QVPh1JJwwwlxIW+IXsD5bzS8l6rO
mQ0tqSRvj2F5TPqX+SzLh7rWRLpxYHa9hj7Vikehpsr8Udxyjd3hzUfhg0jkEzl6o2500gDDFHox
9QogaSdLxavGGWm59HhCaikXG7L/BvLvpxLeVFwIFeMnVanU8ftNVzCJhgCrJd77SpNYJc865rlB
lCLq0gHDNCDp4fQOM1D7+gN5LsOspSR7LsO1jl7ZDWje9gpQBtLx+aLtfXhdZQ1Pv5mYTmn6LeWC
P3a+zx4Rg8VfnV3bxcCWh6w2pVFLyiYMyxRPzlQpa6KcEwWWHT8KmSEfrqdhIBVZuTcmZbNfOOBr
53tcKvAOwSNEQJdazihZ9BM5kJVSI+Ng7SNxKjkiHPs3hmpPZ2bh5eyaiRVcJk3XEbe/FCIjHaFw
YAAh9hwyhLsCkNDERgBjif08ssL6puwsiutrydkVtsR6OwpuReqKkAFqHy3/FaeRuiayBdj2BIic
1bwJdZk7VOSfeXKgUGJbk33T5qFDT6e9crlYyuyxT5CABeAz6rcfht+8N9RGwtzR9hCu9jD2DhNz
v8rww+nVrdcVwyuyUjEtFByuN8K4r3G43246FX6nG0voE6IX9Vc3y6xSrqhWO0pWfouDAAaEAbXv
69qTTSpw+vP3JloNbz+WsqAtkwD0/z7tCiKVCEni+KYoZgTgDks/XBnpWgXQdPnVP3uvDRjSnXB3
C0Fc+AXa3Lkl0WvXsr9hrm6aewIYta0CpOt/xRJe3j6/I+BvUH8ZWGgvPPoDCvlQEDFEQak4siE0
B3cuNqYK/P3YjEe7UAZulSoSDkXN82melx0Dle9UJv4xGwsaFKEyyToIgHy2WxSciAinK0LkuRCH
r9ZCDjqXoOsmGJZ4xb523dHcQRIj7rjFtCWedAjPab27mgppBKmmVkr+raOn1ru39VUhmYqy5j3t
Iy/JtJ+vY4xjcwgQCvf77vLJ06md09hP8qxEjFeD6S7rDScPLYFELw+4bEtcarFlcea4ZgXvZ+vD
97xSQvRXHjBnYKnxvYMRSBQYdQrwBBMIPXAn7gYrad1mH/bJ43r+DTAbYZR03CWbmuUUbQsO5Xc9
inPZGV7ntXgBDYVkCCBiqRkYpVhjayV2H0OztT5zlckY0RnIr43kjLAuhVUxoeJyMp9U9UsGEL4y
avWtCbukIdGHk88TlKm/42wpEHVDWNW2VlyxXPh6bZGaKXlZdxVEQLjNkEv48krk8yQtBXq3VZIJ
6L1h4IPcR+sf10oCgK2JzodCUisbWGC7KDJpXdNNXOaeDUkofsryqJWtssMqF59AdmqE2qNRpWmS
pwErVHkSLfsjuiC6P3QJmt1W4S7Oh1Og1IhkGzSFbxn26D0HEEZkP8hKklqhe+Itm/EhY+QXYucp
BLhLLUyTqCdiL0dwjZNEo+e8iC064j6lxhDo+xw2mkHV5IKu7JuvjTx9yxxFbeEizJWT/bLgOgWH
jV3X41I7MDgvgsaYCeHLPFCXbKw3/+q1O35HbzgvH/lDA/dFC/ZW4b9ggchj9qemrhX55CUS3Xys
LGyzvpnxICC/aGXt23w043Etjp/n0y4seCTZvJAJDG3yaeyDf9wLPEZp6OT6UNPLOCpbl2epVIHs
riis/fNzlsgYcNehCelTOV1Pbnnd8yzZ8WRpdpUcpqfX2DibG8wWtlRHekSlCJfBxfN6hzzHOf3I
uHpWTx1t4e7g70l+SOlZXJFE8qCXUwN0VcE/rXMPLTWrRl2fYCk31X0zrT+04GfyulG0t76uzU50
Blc2gVxaJoW8DPVtOt7NUoZh865kVdIMFLi7+ppcATwvpkOgRRBgVFViDW6FQa/WIJyDgkVmAwID
UiayQFZqzyOEbh9Nao51xr6ydJ3v535YMaL9vRZZTAKlcy7M0q6mo9ELVBd7KEp+dQusEVSTk+gU
CVQVdld+k3hl/gn4HCyOwEi3fxxG+SdygIGvL2rhwHc2GNRSHNmtuoohU35f6R1UnsmdVeQtS8OW
fIPz+Picp6ipRItnqb6Xytxin+LAZY4aRjYRSPHgGSj/IS9u/yz23rhlDo8dW4wPgfUXX3ljwjmd
++m9YNFFgoDb7XWdp2jbait+xfxDxTuxY6qGKW/PaF+U27cavnfNnfzaAXrygclVz/HEx1dvl8ux
kz2LWS45FmhZRModuK1/FSbROkRowhmf6oNd/y+J9+ltBMA/VVhvj/R4dKZbbIm4ivlJxjnOqeeU
/gb1+aVaOCe6gf8RCgagrspzWPsRvrJtBrBxDv1S1LNMs46pZ/ddgcujCAlcsfs8DOmcRNM7Orau
oJ6pcEvgjQN8JG8OkO+7ex3NcJi42RxJ2IMk2u7euwwa6fdp10KSPV3GHcZ+JpHJ4VGL35fsRZ7C
IS6+NHRY549Ln4x//bpMPjAzQ2OdLUDXrfNbrPKWNUan2G58126E1izGQwJoIzjAg4xjnBU1i7G/
POl3Y/3wuKZA7YLgp2k4bZqAdAfDmi5P3EI0L6e9IuGdG/SCacF/S9uXNnhYDqmoSdSYJEwP9lmN
TmzdgRmUbQG7pBSnlamUc05CKW1EklHgLrkXaQjbsXB5oiiasIBiJri5aFbYjaUoKwVN0iY9bq46
HqziWh2qbfLyhPDl452P65jCV6VNWmEHkNc5FCnXCgBiMMRfxP8cpXgN2irLsKgyj0HKhBv/z8oh
1FBhpYhVDs3Eg10/E++VOgpIN3n4fFoxXBsHWVX8RRwrZNxo8XEQsooEzozQhGuqYwD6m5Zp9YAu
SLnPFfv7Y1GNrKiMAbFcuYFMGqGT2OknKLS02d+GrxYriKbh4lbNZ9SQUxvHO5pJQzIb5raYgYVe
tiLwEWbFFHqoEayAW1q7HPIpQzEBFZo2ehmBzAoJEVazmHpL80HP47wdwakn5seY8NNj12K3eQTO
+4Dbo0kUk/uqol+arf3jHbsPnxjOetZMnl0Z3jBKM3nn3SGjSbS7abLMK+HTpWA8kw+sm4eEyeog
nr+IpArxsB9uZwl/RVwIcxrxoHmgLEcfRXFIs13YQGKqXTnqc313QtUM2+Fla1faiUyAbe88k9rJ
1RGEgeBhv7bOSZkZyrAl9dhzH+ODAnJQL7RPu7POsKenVNPAZzhFwqIXtZ+KlwSZ6C0Okzn/LRC3
Mg23wP0EBNWmh2kFez9gd7eZiTkJ1flgEwf5tTPz27t3fMo11pwSMhrQyOkuimQIjnPIbu0/0oFQ
q/tJ2/Zp5xlAKQnlzn6j7Mfj4i8asCkr6gg68Vc0IPSPh/ycsZSOuzdwQx86mZwPUiuQ3Q40eEaU
ZXfr0FfWJsozmKdsd6No2pDiJrT7q7bdmJSZcvfPBlg0OEiOvY0iecsTiYqFRDFWWKoDHx+ZHZhj
WsfvopZm3DKQAeyb9o/613Ny9PmE+Rur/jTKsKXF1zmTK6zwAPmj66SIDtOJC+wiKh3t5MrRba+T
zFHaMb/SaFZnd0piLzXgeZaQOZ/zuXbSkhyYhNWuxFF7SclJnuowIKWo1BYClBeWtLoVWLseRtZ3
BamaQY5R9S4qkcOgeGbTrnRU8qX2lsk2BM/GSeAke6MePmkMzOYSGnFstnBPVE/J3cAVUCkuQ6cR
6FdGmvYs9r6N+y4heqInobv9LJh6u4t4VtAL+taqtgaoFnfPJr+aFlUd6w3PJjaojeQJUg6jpsMT
WP5Cx/WARuvx+gwMaFmpiZu+4bsjJcEBg7IN59o90c+8CIn4IZfnXkDcHuHTgfNkHtS/GEeqQ3Gc
2OynNic/Fpp0PoweXbP1aBkaJx9GtaBnWN5hNi1NTm5zkaetsUhczyFZElbkCW/a80VQOjyDSlUx
lI92S7hbthgfN2Ob+GfFnfZeGLRsBrlVZgZ/lobr3A1mnFxPamyiGKc2Ig3RGi41ZNSQRBcA++he
AwSic11d6ycoTbYoK2F+ixfq6rRziRRLyxxYkfDGq6O5jkG1nfPHjjNKKbZkRENMEGHLD6Y5C22G
ICusK9sWm6I5p4GSXAzLCswSsTIjByivx26VT/l5ZMkx/eNeC/l7DKKRmgfPf5CgoM9Zy7TSQ68K
/t3+OqWnUjs0FyXB8q61csfcQUWRCsq/+dgCT8pOdU2qaSBcKVrC6YjNlzzlOYGGUROcQe3N4m9v
/OaXzw5cw3c81Xh3h+lW7IO/01zbikpXc8u0O4OWTjz4YRqkxMr78EVtE213cAQtIgb6/OMjruQP
Qk70zEI2mL9Y5bEnScx+VGy5ybf2I+OfPSGgMyxkjqnwPourKDvDqTXHN7qlMgTHGNjc7CfYmUf+
KCRQ7dRDMs4iJqsyQFuZnemRy/SSdRMQdR9KEd7KCryEA7c8GwgiRQy+FC3iSHelPdaFomrdjspp
Go8RD+jY0fjaZI3pSLD6cnIgPa/3NaU1g+KG7r5r79/bxA2ii+baNPukroU8tjo1mHHCIx5sj1lE
FxVIih27yO28YyXO+kHTauaR8qAlBQt+ly/TXSiCP/BSzoHweTsz005LueMHMGxB6vGqWHbDKyWg
uLTEP06U7D3N6l0z/lOiPalxWZHDZwml8fY/ciXLPgZ87hGHtHJV/FvJ17/d8C4ue5b43o9bOuaE
qIwsMt3svUPoNfnYlyqrkd/OFhPdHNHGwyLLi645qkGh97TYsqpQ91qTSLMebaG8GExb6wXcN7Em
7rpPMH8LXu+ZeetPFmLui1QEHFdg6hI3TPIqIu8fYdG475Ie8I5mSCIp3okuKSpKSve07BcYE767
h60I7pbxs08iSCkDg2vJYhMXg6+9drSwda+jJinBIpzfZpr/lCjqQMzZe6+j55twbsLsAXXVKVW5
S31k4/hjANnAUAIYVQ9Ht/jL61ocSBfDo3s+nCeFqQzc3wDFHfmIY4lzZQr+nJ/93YGXUSPbyUDu
cf0TU7V0VoFS8jXCpTZqhE+uRUPKkwyLfLVhI8CTHNL1PbiTxZihXFqm5sAXGgLJ5C2WTDug6bwh
NMsesVps3exDmhYlDYinUXS/rfBl87uFA29rRLOe3r1C7jV2ce+jfZHiqP4vFGHBPETRh9uBGBu2
6atfwF28a8Y7hWxYpWEHzr5lnwr7SKjqKxszJat3jR1OALYrMjQtc8inxHkKnhWEpfKiR/4WCTgQ
LqjS2Ltp/5Dv459ETI7kOdwp87z+OnsbJsXE1tTycHENrVSAojfMiNJolj+Ltw9F7Je+J1+p6kuR
ZcEf2DikBvKzXmNOkjNvBS8NtkFPWj+7x0esN7og9LbNpGyXKdTdtYdcYkpha28CbBRQNwlE+HGn
ZRxbS2JPaU6NdUl2ZK0ZlOE01sDeDYoR4ScEqmUNLhYQW4nwqJXJaBQY9sFPYQ7td0EOyXJK1dfB
SYGVC/xcR36uXDf70cpusCJbN9O/QTbpddd5q+aZcBikvffzGOaIDQBl6juhwHRtPBieYkJIntDw
j5TMpyXfgAcMubbpILhUQNNf19wTs4DTNHL0drodCyeMYp8sb9t7ePJ743NqAGnJ9n3uwN7xoGpJ
L42826vrbsSJBn/0eYG2xrV+xjgtr5O6XxSMD3fASBKO5CD6L+gjwinJ/5h4dVHJxVRyEBx+/9cD
HQIBtcW1cNONqEDJ6i3ao99uqxyJNf+QVBi4DyWuhK0bQEfeSQhEQyNtFdMMWvbkj+coL9OREIml
RTyaywOb36yNAAXUJ+CE8aI1NPW6pzEvybj4ma2n3MPhbDsSg5B8iZdB/+OHsDgRG1FHaIZGPVW1
AKCZ+zksPwFvaBkT9EwDEXwwkM0rTB5u9LDnY3cuSnDlxwiQlzXZZUjxNmqndwqrgUua+R4DDwYv
PZw6qlceSFaKYtfvL6uogohMuXnyoWSCmKrbnRTeTGmHnBDSXKFWHUQIiy4CPDYF43DhlcNaZ3Ab
GPBfUkuJDXzwfRAMAjiIjLEUqLCVd8poORWfKv3jDsZpQqtNxg4lwYXi6QUwkwdBvMlQ5alWiTOr
7prF6oaYk7tnfS0R61ESClBLMasuRrRWkdVXH8D1Fi+zKgFvYrIvWiN90xFKNDdxLzQX29aDtTsY
0MZbPhTsZ5srR3u4fYsXRb5i/zzUeWFpnQkkF/WVhlHZD4kpKb7oDR0Z+ybeeZG+So7PvF4P3yWd
4iBHDIaW8C3RaAG3pEv4Wm0lbHMyLIDkLZy41zFS+weMeM8K0UOZAnjNSgzsaMbz5OBBYHEXC4lj
Icfy6uKcXNZ6n5egVYo4grivMn76sD7jDIjmN9n2fRedRkA/0FS6lbrn7fe+wBVBtTK0rZuDUgQf
TgZHPPwTOZ7puWRs23w8Rh9yVNYYsV6EjI+KEHuGlUlK8S+JzW/ClDPODtIoXN5UTEcVJWxjIJsW
yITx9MA44W37IcMjmqhTzYJ65tgZTfGg8tqcIgxfzwR4h3gGFzUmqlzntsTChNbO5Z/vvh+T+RJj
JD9HDeq+rFnvGn56tROWGU5a4AlZk+3JwVVDElsFWv4gqO1iya53t8HDQV9ugIj1VQ9P6NeFBE3b
y3teGZWwwSy/f1DW3Whxsnh50Z0zxikuWsd6ou+qR+LctDLQN2aYo3W+xpbEQWlebU6P6L8NOFlH
UiOMWXO3HbA1QyOU+OsN4CE1qpY60RWr8EZyBZNw2v3s7FsNDhrsysU9pxswKAVve9Ufc0ALiThR
xU9EtmXY7m8ITUYi36LpM//DVy7S2LEVaXsL2yMPbvKkWkem7mI4KI5PkjviHdQ4eZ/sZhprmObr
Wl0NozewY4mE21WUt7hEA2ZoSKUzJmY7PHikm4pnFTl6lKXWCuxWYy785dt3qRXwFFt6U0eV//S6
xZS5BQ7Fp/syKLhBbkbKl9RMuPGSis0v/itvL/KHvZarvfUVKr8uDT+Kc1L/zzp1wIhdOUe3dSO8
E2BrO2anIlwDQ9eHsPICZnShBTM5EoHow+OCxnHFUx/4cCoN2+jmQGfLLd/FrDfEtcnTK4XXd8hB
667fj5rj9vQvC+UJ1sdJwoS2U8s4myw9gs4pRdNw/hIrJW4UAa3+nNnRhZCzkJdjSNcabqdY3SRC
WQkPLBubni66ZlRPfN5G5PIVjayIaXVNWEC+ZeLtRLClFeKcA4gEKVccz6O5fm4TPQA6X77R5pmQ
R35x1kJflF5QNFOoyIpnnZ3A9RcWk9k/g8awHCSEWv0k4k9xRFvfgC9nu7R0lQy92gXY+b/KVtvS
RRxH0x5I0m8pPDQJ6LwwY2eeiR8Q6bONpYPLHqiOB3EY8Q6HKC1o+nTKY+1akvhMz+jvg0DPXc1q
Sx99oBhvVH2QqIBKZY34a5hw5VAKUR1nCO+lrpNY2o2yzI34SPWDia7379qDjNwvjLIplsbzRcDS
1MFn+lnlYg/0OeagKw4r3Ya7b64ZoNIZjuDlUlZ79Ji9Wh3OFRBgqpkOMz/YUuwY2KSp/hYw05UN
VOqBYc87GuKKmIinY1XEB6mSD6yhE7ZRFaNL1vFTkjqR7lEXEY7o34sDUtuoh/tkeBtdmoLpoJuO
JSF9YislmhdtggWgJqO2BNEphCUJWt/dQLowuCJLOT7P1R0WPWDOxDSoCWXZi1tziZaHYobCUFLe
G6iozQ4x4CI2tMz4xelwIv4hB889zKOTQb0ssyIiwltIQb689OxlAOW/gm8iBkAkvxtTf23S4JGs
nFrGBvDfBJU3QwavaAn8Wa9MrDBjXrcB9/PufwqtBpzf1qQSdM3G2HUkxMUSDyqmwVLa76hzDCuP
eX9mvY7kOD3qx6uSzUSLCZxOlX2H5NapLGRzSN+xv3QmZsW/AkY5QSMg6q3mjgcXPPADVTM8ZqAS
B01xkSZ36vxGsaB8jIQiJbTvoxJSRjQSByFxsMyt7vKCdvZsA2czcchmk5eZyY2p2jloiXktI6Zg
zz0dyxQLWrMJzfnCTMG1KBC2OrkbQisMAlCU2bApB5QY270e06Xw1VnC3xpQ+Dqd5momJT5S/6Jx
2vtKNRwDzKNrhbjVXWYFXhF6ew4coNAA/yaFEjZ1MQJ5DEoDJ2ejhUZQoMWMLujeQ0tYCRHris7E
ImQgGhajBoLuD2AFWlDcOzlFPdvcYHBgT8xDqCClKOJBW7CnousRLB/wYYd9l6w2c4sKQ01Usb+q
+WuefL30KdCOuvyB++hGJ/etMkQBwRlVg2pwc0HcCGnS9hKbLYwMc05Ii0jLtGZ4Dn+yhU9ZZruh
uq/5THttfl5NaFvayNOi01KPNL3Wsv+3y6cO96GJemN/nGMIkOGKadW68H1nRFkvOuMkBubrcJDI
Vqjs8f8snsbZeL2ZEEnnmWZw1Y4zHbK85shIQcESHj84yzRA1S80/OICLoD9UG08Sm3uuo2Fxkpw
qixcggsybLz2akLADUXP6t1uXs5yQCjlzUEWhouryPasSbUV9RpGGDQ5m/Qadq2yZ8B7d+23HTie
U1CiUgt0ZfeddS8rMKezQugOc9ZCOxTKwkYah1M2jYU8QIU4+IJzavxQrr7C5xByaMYK3t/d/xPn
Uy3cGj7VO40hT+1EIyEnEUve4mi4zyhYFR6ZUXjY6xWoiLaRibK0KvMQV5C8bup/b4ydprEZjKuD
yejLo7hwyTlZf6HECyv9g6DojWspufSdeAuvaXP+klQ8Y0vFvpS3U5gaVxqRLmllHIrU4Z7tHNt+
nrkMtCXo33cyws1ekVcLDGVT9wX4Q1aLcaXVWGM/0LKX7vVAOlc/NOTvJ0FxzzA6ODzIMI1tUuAB
SAchw8B1dMoyjDZIuqAB6LHDAOzT7D8I0PyApMDraODGABReZsi5wvyiZaQCTdfyi3mfhiqut+Qi
GoYbP4HLrK1K4YiU3EpDvuxIJNtS5mnV6CePVKJ3ljzxNo0ND6gLLgcJM7BDRlW40WORXVf+y7VR
c7mIKnK4g1RAGqV9AfqMG9uFQiGp1sIURlbkZNy721gdiXxYn15SRyJHzklYC62JLD3wE1KTp44v
v7X1IB+OOKmlJVQuVlnE5VDXglov1Vx3WN1RLhcRxBfUzbOY0w8hEtJLHfbqaOeQog9K/I8L7gT7
1SoNDhDXwUkF38jlqF9W6WaHbOYgHX37Yu/pwbPc7IEjG6tN4q2fdYv/COqBP9alaxBMJlAEVxY4
d3EMeRBBiZQOhrsB43h1cwuXX6Rj5dZGH3l97KS+Sssz0olHJBla4ESUqqzKM3GZ9PrvPzDc6Tq4
ac5m4UpG9pYM+9SmZS3m3bgpDleR38PqaAQFb8vxyydSlOSsVwkVYEqSjlYO1yDFtY039SROfzNq
vhl12ovxhXpyVjiZv9tOoeB/Od/ekUUqb5j0kYkYvL3VlAyWxm3VjgvX5kH98ud0hVGt+joMjDKZ
bGfFCDPkmrUkJSPbf7WhrTYs6LTFQ40C+NhE+e1/CG6ufbUhIiu2EJ0AFYq3kOeCOztSjMyhW6Jt
wPLCvjBhWEGCZnZGbdCD2uFKrbUV0sMacxI2SWgFcYgjuno8MyzBnejkgAtzj8olFYPJc8zN6ARq
UE7SbQYfIMlRBy9fv21Dt263qxM5PiPkZ/ZYwux4BcWjQhAC809+fW1uV0y9kEeGr+hXd1N6G/zp
AhDLOrzeHgCXLk1bmgrhxUXdFtn25xDJW3fR9ZuUk5DHaEYcsnDjcqIKxwwSF777I8MFmy4ag4F1
iAZ93uqZXB2GDbCUuDfIzmu8n+m9M/BGDXJSY9DYtG9FQP1BT315TJHCPDIEoXGOW1WbJdLny/a7
mAUyzqVylP//MLnvN8xfF2tZ8RfKl2PtVMbiGd1w/P/gHTTEfRcAkv0CnUyN9iz1wZ4E/4Unvr5p
O0wMx7DfY26fZJXEzMK8tFKS4z3Ms/qQsRpiJ25NQ1GvnO4QsTmQw/VU6Cn4ApLYBLxrK+JxEt1B
3KHx7Kf9aCSf1in0YWU00WBQaxT3uG0UrukDOJG6W54Ug4O92/PbWCiuhyUBZueuVg2W9kj8klYW
v9cu+yYeSySWcx0fDG+f3KxvDXvQbSrVkY5q57rD7L9QayYUnmEwaHiMohcI2DaMkdnHGC62/CWF
0zpVOJXyPy3zLJUJKvOq5iwglIq3CrcMiqavjAG9u9q2EsHR7odTsiqGX7yUrVfJY6uTjPBSA9N3
/QbMQ3yRwQtenAbAWJ/TK7zfZK572EH/pMMq/yCOGWsMV83Ojs3MSUGgzy+Jv833Xzcp45cIPOsB
oSULXjBAGI5bzvO5r714ayWpn9t1FxQo0izPUxuluB0cGmTGpgcq30l5OMK3vACJg7upTpCm6Fp5
fgYr+oO/mGD2tnckHlc4Sw5klEaWQuCR/e+yj8B6lbtnReVsW9S02Ewk0UQPri/qHSqNT+hk92g6
FW6TY+xAD1OH1eGr1xh4Ag2bwQYEoDY+sNWBaIumM8FBolimOUBQxMcUD/vPaAvXkApwFIJJye+j
S2W+NRSsZJikAAcErfFkUTsA9cTeuSNuSA0DVcvNkqbjQnIbYqor7TXMHGm3oh/Di1V7K/mWNpgx
0UCbTr1eOOw+C4c9q7sYC+qKgzawGQBw/Yg2kY1IkB7Qk9w4vMxaHsYd9TCMde8c3qisaTL2L2H4
XqcGbXXniR+kDO9njhzBVaex+tqN9ZrHHvTV4ZCDJHorXYZPA2+a+YGlg3wAJbbXUoj0S4swFPKS
UR1VCj79Z3O8EpxTtGZ/20PjqwcY3b6mlh1f1NFFO0q0UoJWTdEe7tgbdd6EoT5I2wO7L6Xmblmj
ALs5NRK7Vhjdh8+JYwPWTa6jakZHdDtDLIN2DfMru79oIdQUmW9wcPQvq2HDk0d09dZFpLD9j87l
K4SFpT+mbZbpL7S8O91xyMgPA/lDKsDuWaZK6kA0T/nNGo1bhGBi1BHy7Gn8xvcRyb7WcQ0v5Qcj
7yasV4EG105C0XDt0E6FuOqYCl+W7N0Any5Uy4HyeSlk7u+LFPMHfMiDA/jWA/40yQzmX4T5NwTI
MT8BmRkOm+NfIABF+IhRPpa5sAqSlaerKcgVjats3J5cW8Xcrn5dQanE4cmFMqqh5J/BKmm2Qu3P
XrwzK/37x8kekZvOA6K8Xq0Q0QjGrFnS/mcLkMUT1AAYP6DGopgbM1pjLIdo9UTXfGuTPsTXamMp
fCh2+mewH6Q0hJjKYsAIg5/IyCuX8dAQddK+llxvHFka9j4sUlWJMDyQWiDLwlDRaQHM0w42ZBKj
VaKZ2/oL4Y3wYGfYLqVxpNpFAuXv1ew2bhqmqBcNu+hxz7nzY2t7DbD04pPcHgVrEZlBWqGDWiyB
NtbRcGi9WnF9D8w9CeGuL51/hcLPVOzgKye6v+j4AlCzQn3D4JMQHeInnXAIW7+PNx9+D1wVxCxs
7nozxIKwX7hSUIyiKaImyOUA+L+nof2jqIFhRdx3MwufG8mJf01ECQ78wq6gBCRlJIN+A9ED6Sko
+nHW1hAyAEMztrdHUZN1dbFy4SAIC2Gb0NDJMyCd24C9nsAnpKFb4LloqVhp0qYaNyK9JrovxnGS
M3tKD68D2zkMR4FvJiVeQsob/BWyqk6XeSfFVUUFHAk+YFRmfHNyWlJ2oSUs4NHqLaXk+UAu6uvB
9Z7jZ/0r9/vRFwDldfHSnAH/vYj/VjuAVwhokWJmBq9AasKLu/mB80vEpCnqWMtVbAto8xgcgrhW
M4fpyCKVkM9HKGRKvf+GKV4PeRnb71xz1jQiXpVkM1sMICR8GgLBNhMCLPmwPcdSLcZX0wdXKraC
BJ7rRkrUtKjAZAsMEGZw5+t05iHQ16pQrYzBRZf79LT7DCyoVArtqq7lZrCFv8n8J9AfU9k3+GRf
qordNfpBQtOp71ZBaHJvYGqboPtjd5kYVCvfIak3RZ3X9Bg6aEZQP2VJo0FPCV6O6O9o8arirZvM
0IduEhBSmRQxJWJhGbr+8S+l46Tf4ctgIOI72UENw6kWbKUVIlZg4ckRd4sFhS9RFurqu7jLrXN5
5G208vscy4sBKT7TEXipCJb5UYvZLflDqLImKJhRsK4X//ynrMc+u74CnAXvCniyljfCgzosHBQF
xfx8hMY4n3bdYYeW4Y894rudVAieBZluNlzR5KRPL1Az2H4hoWJzqdiHbyTUhXjEDwLW6NAvI+NR
gH4Ma5i68wYF1bmOsQ83ev7WEslxx6/Sr5OC313r6VM1aP804TWd1dPTozoXZJSwmiskIIM+3/im
SmGBZnpL3txfb4ZQx6xF8/GtjdG0lqqUl51S3n7p+FzaasA5QzjCapkQMc8vVv1sMyTdgs0Jz0J4
LFU6xwrpm/NLQf39xCiVvoYhU+fxUGa3hfWkl8jmQ9sC047RJ7wnUsNoudRiLskZHavOyQ6KGAhm
7S2Jma5b+xIitkuCFGGR72+Jt05nE8hqZtXGZwxtNqzVX9r5YSIuLqWIpvjWXci0iHigEbGbi9Ae
TRpMBdqDmKCQvUBqWuelchPa6QQifilk+Akbs/jDAUYOw4Utu0YFbb8+aIP0XN6+Ixg0Qj0duuJ9
p7vGH79v0/7m7jG3ZckEETN8I4ODDuYfmbeuX1lWYYj9upvmC8b/9GmjyigLr8y8oPViW+B7XOWW
npCx+obJ8FfwDEtpduJiOPM/B9Wtf0XUpTaSrNlIi5xtI+XmWQjlvQXLuWkgkICIYW3G2we35AW5
KIH6mIGBehbXBpE66N6Hjt9Y+M4Fsy0cD/KWBgywTbtvQj+fmAoWxhweFSLSi3yNyiNZSldjzwea
lsZP9GT8s+FuMBeK9PLAd9z6QCVkIjG94U5BVYyB1HznJsP86IP7qftgrrMbF2VZtUwZ8mWeGDn7
v94ccnpoGwjCsErtY+Gc8zyG/WVGRTtBsRD8HVfIwco9Ngagq1c90UDLxV6249F1S6u+d0/IP2QV
cH76MEPt0OwuOdPvj+zkMRiWbpapLFwFmYOzWJNFmJmIUfIbd6uZ7ug/n+FDB0BtZT7cCFgSBzem
QmCol2yEHgssy8SY1a6MYiogrol9Fa2yyOJOAwsImzB5lKYi6MDlgk6FZfvij0wukKfTfNaF+vqI
vn84BejsP7prgi9Io2OumiTKKfwIuCEMmv3s/eJY5oB3+1Ip9q7vr+CRJ4w+h4NGgxayPLm0lHGE
p8GUfLAPCri98PFZXEgH0l/RV4rFJMi6VhtZcwC0WhyAllY4lsqVzAaoN6VBCuspSNLQBnRBmCcW
o/yAiMfDkeTXv6icHTYlTjJfQqgxpqLrsAJONfbf1v3iXHliiF5vJgEl7ehOUj27i2IC4xBDsX71
vzCUsJDURh837SfCx4IjReQ6fVb2YJv5C7/4M+0sAWryZitqL/VEIoszb2wjczdplFTjDvkj3vh6
rWA2VdfBbKDAmycgMScsTPuKw5pKNm+XLMFb4bgqxkOEVH8DxNpoXF3/IpnihHe4dBX4NAKQ+oeK
IT6K0g7zrkabkcYRgDWxSEq47tfnOXEaPTq6maxykZHEFHje6HCE46hhSSenXnlzI5fbB9YPyyC9
n7ZF36u0rrWPCHIkzV7CGSb1OM27uak22PFh0lzYqT2b3YlJMbd28qSiQgdC8/uaOGPkCTAK7Gs7
qU5AiL3+kNPkx0EB7oTjt6bw4etyAYt6TG66Z0iFRN10/rTtDwP4jYMMceh33+aisn5cCa77Ns46
pNygH5U/qm7sljoDVTpoTJr7b7WiXWz4MXp7uT5sfko2PY4q2kx/lBPpArCrCIWOpVGxbw7dj6OL
LzHbkPmFrgH3nsc2sA+W1CCm7U/PbBxti1MF2ktAsCwPsdheOcvQ1OQajlwv8Oqzff3lDmiLSYnQ
3OANQSwAmRoc2bMPDxUjiVwqBv5BnE1NvlIb+HUsG5ISrRVYr1aaxYNPIID68yReRIsQZpPTcCLF
mDGx+V1w+HNPqV+akHiLGY+wp7bnbdxZ//5wlbo5H+sXmVCNpFZ/6hwDKM/d/t29cuHLOwSuJ0MY
IXSkKZKkqLpsoaMNCCpnNE8gvelcG4AB511pawdSzs9JBzGAxhBcolnLUZxMevyXwZPh1dP5SnOU
v0r5RzkczlKbt0Nsxu1oMGynragQeu7auzrmEqVkMYOl5qI36QSFpze2/Mk9vzayH2Ie3z+RP0BB
e6ULPAnAe4DGLiGNbaelJPgaPPdxEM7H4X9Lx2wUMRCjN3fx8I9ZXEvpc4SRk1JVhlGMRVN6WHMl
c6Kz4ahWH7kVfc2ZiMsIlG7HKblfyRtnw6Xro2OPWuEW1aU30vMWzCuprg3oyA/Un887Bhn2IZ2T
Ic99KMU/JINwi9w6FMBzSbex+/MR8LXQrgcdzLAZueYo7Ljs5GwehhFXSilfdK+meSQxauKJlRZt
LxKu5FsY8S+YnlN5JrBxXZKsTmQLqrq+N9rwYUvviZCylNlI/ZPfsm/sRUIrf2hcEcn2sk9+DWxB
+PURQ0AAXhZrx1UmJBZQ0hPIVpXKMYMHE2ICfV2YsN5fMkOoRnUIMt4CHuC2bd3tt/iClkfvABxt
V4EOt/uzuAGybtLVsBNOyVuGikKBF8c40DCzOjsHNWCOiQwmmt8Dm6dZflyKZEms94N/zz3e1TfO
7vfDMIZan1zJEmpwBkqzrUWWDH0ONN5U4q/Q1/ehwDdQRPmONYCT0grV37VJCsBtcl+xa4TQ6LnU
ctjwDIBct3t+0MQrZARSbESSrHNYvhUvDvT+y6BJ/sycRa7aE3FKgH/OBN/suvCiqJQgwNR/VPak
4lpi5YoOHJrlnQ0TgSmDPjS8JM5IhvddtRZqfXwZ+QV2vHyskkXrHDFMDfnxeysDvKRPRZ8UsB6j
KDvu3u6TMrsQnlkWFLJX+9RreAfQaB9R47BX+vsLK9YjkSVstW912U5kVJxWbK3PQv+nOuJvZsMC
zLZcMvSNF1Ni/nvbyTkvEEBK8oyqg+v9lTZTu+VSMiUgVtfYZiM0VnFrW3Ii8+/fhxJ1DBijqn9/
ZQ0RGQXQn0QMoSV+hHt/AWIdb/+G2iyWt2p9qLKwMLey3fhZFYQPxiNdcaVscVmBLT+nFNef+dTL
XkX3+vbdwv6IUCBXyYkEkTusgSMPIQGoWjMIDSbbmR4AWjaq7HsdrFc1vlWQgBw5M+fY6OJnvZTz
+FXXJXMj3SF5ogTazXiORdglgJF4PmkV5NCXVwfyOb45gdfX3gpE/L9JJR4YqinetphKpFSVQ1AW
aImDVCyq3YLZwY95t9WW9sfh7RGe1oj/hZYg8hXhK5YhUrQxhmCchJzz4qvcWrVLXm6zkK0j3XFd
lxRsUscm14ILNgaaDEs2qO/VzQMx6epsNT8QLvJqq+gVdKc9DCGDW3kDzehi6oK/LM7C5h1ENZ3l
mO6WwUIrHAsqS2wGGsDHXebvEt+Q0dxmInn/1169oa1mIVbiYc+PWacbIUDuaGix3qDVxM7kah1O
sTpZ1h0Gbtdzrb7V96HmA329chlQcZDK8//50iCWXa18NTGnMWf8OoKzMsgv+cIsD/1yZiZ8f14R
8jgfgTSw5/0HucZaZm6MrnFHX471ZN8bUAuZXqdn2AF1mm8x+rlOMjOcy8Zv9G+t5+dVl+GdmPuv
Mj5ko/FMaSSQjl0EAv9M3dkYnVSPgZA2Vix5R65gGyFQWHcq7PWydQW/DPB0IgFGTcwm4eZGcohA
jBP4T6iPieWRFbjIyu+g71YjWC63y1Nkd3hSFEek7nn0u5YhWggmL4bIwksdJSNw5SdBvj1V8E1s
UWRpTlPp+KdQa6HnhGy2tTWzmU0jwSSyMkbMJsmsz13ekf2z+oFR6YVfP+SdI+0xo35RlJf4/+SF
elKL+djzGFD6wG4tqHhk7uBBm14tv+xIvCHP0WtIAMHHIZDwRb8GTcx7oae5qxmkPdj09ADKeQLE
nUbuTqRWA5a0M8GImCAl3ApDi5AZBJRDKubuhqfZIGZWYmy8K28WtmxXZkOYPvlExkW+uJpTO1W/
eBMbPROPMBNwJ6Muw8mSj+s7LKMKI+iayAQf41L1A8DlTrnE1hHaFom8f7oTIVe0YwTZjWqEm96j
fHAU6iVG9lkzmBQk1PQF9GhVmIR0h1Rr0LRc/Z+xeXCVGg2Nqiz1cxb3ec3ATImJukj7Y3X7sIgQ
IQ6LUxkKoJ/Lj2URggFPfAEGqJsKmx6jKjQCg8DwtkRb2lkIPuosByRnrjUFUwDA73Q6XZasMcv2
hSfp9idH+o54kVARdCPoE/h/ty8yzvJ2y1UXToVocyX+HN6mDKkvgwQDKweIyReoOQ5GUWBkuIBL
tB7DMWoX6reJ999TuSY/avuIxh59G63sPUT3VVSHu0LOgGIr6zZd6R8IaQDsZz9BCv3J4/GoRsN3
y73FHRGLWunEV3BNWUJjYN3WTqJFN0IYTdrAZkmfDZRBkVkWQIv3rQYxLTYfiZbZurynDaIjAEP2
13KjgXn07zZNzO8kvvuwB2OMRsRlbn0kCJFvxFM9PPPGnvRm8VkPQhPiOO+jMc8OxmxFsZTUwtk3
Foi8Bu5h4UjiraabiBWZh2MwJPMGI/SuIHqoz+GUNFTxo1AC4H0YZeL9R9D/A6EfnvS94OmYSQ6d
xAvDDq/KkE5LXa2QRsLFgRUECh53eYSC8ZYr7PU8KmPXfTx0fSP0dwLYomQADlmMFzevKojr5Js6
HRRJP7XsJNJ2UNJ4YUqRQz7p1evouSUvlWcnF86lNuqJUxG6elK4YBChxQ7skoSq3PbKqlJyl9WL
o1uKk8beCwO3Ac9b8ju9W0PeK1YLc9YI94fkVbHYyDds9k8zIGbxp73sEJgmwBIrVHALK5P9Z05M
yv3H69m93Ck0DWnORjuynQ57zNqA0OXekAZQeYGAkhmANdqCIzOl17lMgChypG4b+k+tuSxFEY4B
mHMD9SyI12Qq5N//lk8mH2W1o2dOezUMgIdEC+qIvWON2ayF4P28eMlW7Wudp9bBZa0oKjcUgwQI
L0H+5AWU6ubE/+mkrLY8QNrP4TFqJLkuLo8WGm/MdfrjKC+d32/W3kBoas1iMsIaeg6SxGgAg1tz
S9yUcgNe8z9wFM/fxLjtjONd/ZCkWWfKUt1Hmz8SdcGS61e/u3dLTJh04KqJL4lz3AkrA2VNR1mZ
vaRTLer0jAC2wUhhDMiYE/VtT/2SI8cA7cus2A4ATDVDYokTj1KfFyKWWUPjvyGoRGze7CIcWClH
J8L6VEqjleWwnSQZv9Um7Pv7CN6heUwztu70+noAB+D/WsQ8sHNVUKDIURyQA+6r2kb/CF4bBz2g
dvOZPuYfEG1MqrubKuet0rmZqYCsgnISD114+IwOMV5oPw1RmIwiO58UfDdevgm1fyNhycn+GiIW
joIsZAvDSKTECaay1f0vYvocI44J1vPE1TxjbUR5N7wIgFbt90BEqyxqIsLn0Ub3C4ZoFOf3qaUN
QOeIbvn6zEeg4+NtKIyzxs85lQI++CVunUsmuX47aC6ysszexPb7nLkZhbPYEKngNdqdkQj1fNNe
KpBQsF2bn0gFMgCiNDiIq3t0zRJMuE4Gy6F/lDWhBMoz9waHCwX47nYLpjkaGbnJiZszNFRPzw2/
2EuiVjmM2K9QhpFtaR4+3+tXdHmGQnbyS88tGqttRhDEjpXUXjThiENWx+KJUMel3J69X8FL4H/q
LJ0LhdM9JFDOkSvuhpj5ATGUingbVvUQ34t4v9dm8WmXU1oOIl+XxmjUKFWZeSuO/UQPtANS3sVC
ZYj45UsDtjBLkM9XVZPY/0hg7t9onIr9qs+u5W2DqlVC0XXv8d5etM8PLV2bXdlLHk3xqHzbGCnN
LkMrB+gmSQCQdp7oiRxQ4EtEFRj+yMjIIOiTy07Fi08bui4If7oTe+ch8ZpDE6f0smMyJWjlrazo
3eTbKcYl8U5BvSYDqhkgJ3e0AsM7CoW837jIIIkvaBFhKGX4ML/sD2aGt6G/Oc2fHGj4HfHqb7Vh
2y0Y0b3NsvAwY7Jeap2/2YfK9mx+V8KRkl/YkCxbaDSseoXzMNTnhcY8x4J698m4ykaXeRfqQ0Gd
7ZOAY91R9hwphbfOLNQtQ6AuGCHOeLh3d9dZR9PThfc0mCaOQZ3QZSgmOE1b3Rcrtwoh3LKYCj4K
ta0HF++Z+gEZrQ5mf6WNcGFM7OJ4oiWKLMHrkj0IBF0aS2K5J9KSy5aiJyrNPMOHebExaaxPH4jq
/zqtLR+CMgeZV35nEZy+oEvH0KT56bSckkc0mixVWpOQihE4WVWnvmdH2PHQmD302aaN+ZOCiMRS
NdqCTJk96nv75ZkmDagBr685v0c+KOJ3Id8+9q+goSvaXw4+ICk8oOyluONGKWyaVjwV/U6HooLZ
dL3prThZYh+LkYIiMpJEKADNuihKJnbjkvI95o6mfnrb29U0HeI2dAPoDEi28rXX3y5mI1kaNYxM
ibFO4ykICiiWJgssQWbotYuPxD0lhlvnOthKMPKEi6o4jvldLUQzU4QFKzqpPhPN9NWciXAP/ela
oMLEK7E4PllnCAq1Q7tyGOAy+2icE2vrRZ4Q7o5PpLjRzOaLv3lnIyrx6WsQYGa6LifCNl4Pd8B2
2VdEtINpbtjftXhI7rj2plRmsGA0Xv9jlBbXUrb3FVEr+A8nwyJ3BfmF27xDDoylTrqC86jnmcMp
rrhAWqWRVVn5+3xIS8W3TIAJti6Mr4LZaXzo116Nhz0LvZVyjFbWRF8tf47lfDkVI4SxbX/PrkbQ
GWcUZJ45BvnIYQFKFwecv2pqiO4RdSDenvM8QuGjIToU0T8yVRSgXdflI6LZPTa16kqf9z2Bv7et
FpXfvSInGR1rMhL7MiAeLV/na1A+64u8mPOJlGtXk9rzl0Y1HKfsXIsYEqG7uac4dMmv2KpzmqLZ
HlIHjnDe6FOCp1h9r82ZfNcpwTLAvx0cPMg7zJNg37NQDnMjMu3FwmER925Wfv70P4VGbEqS+hD7
TxsG+43b8+up5XQd7T3DJtBGqd329aZo6HXJ2itgoLpHRGEjJDxVqRsF74XP/1JDfe84R/0TzD+l
YluGWsjnVyJz0BdMYdvMF06Ha0GsWzKLM4eaW5eO8RokgXtH+5RIt2eGpEsw0hw+75+2shcVUOC1
lBTvKXZ5ko5Z2qYHajsqmd311+NbPQCEnRYXKhuktJIfNKCQGBuNez1S3JLUkpZC2LU8fdde5oUO
2sKHccrc0J0XsgzaMedy4vgoWaoSxz3dApw8wqcfZgJRbw0ucKb/r5S1pMf23p1+qHH/WVG8/1N6
YyKLU0UJTZ1KEd3YGLrScnbnSY00EIEG68y5Gy+jTqJL8w8LAJFrAgj5zcVqhylDVU8ffvrDS1kA
Djy8qNv9bMUQVs25sE6Z8GPT0o1ZlwauItgLGb5KxAPfmp8nJxv9L+FyhhIbts/LdnpC4qmTZEU/
oUQPVmi5gUHSfdQXa8SdvlBvhYv1vO0XYDc/dlCn6WZaGRkrBjmnEF9p+RNllfWAG2p0nfwco5PV
LrUGKjWALFtT15pqKR7H8MKP+s0xhXhx/4JZ74QrQZNjjtWWChslGsqLU4JgmzhqPwIXlPOqG5xN
0W3bRiAXzVg9VDU4NBeYxWk07zU2FRRNb+Luf5ypkri0cGkSw9th9ZOn30WLwoVfTPNvkuZXJzIy
dqqwzElvRkNm1sXNNykEAhzAi7AZaHQkSef+jNn4zSMf2+AZVZE9YgsHIz0UidAJ6FwYb+gmRR9n
ODPCWx1iboNGylRd7kehl1I/VzSB/I8frF4bs9eFEhkmUjeIHwMHPvjte6tBg+jtpaPVSRNXQREW
gy8f0ZfO45Wu4tuOj3IGmIEJz1aMGXhDdKPhhwoM+M8pegQcWK6C+atUz4yAFWZErrLSjMhvAtNH
K11veJdOOFrOoE7emfa43RvI3fc+1oydSsnOH2lAvwm/R1ywa/WZaURn8zr/gBJRF6nd5mUqyjhk
2kTEvY0J3mUmG7XCLoI/Gl6Nt6u29RN9hrfd4HwAI+M4XAKyM+6yrm91GQq6VeCBEIHXMgZ2mpa/
iUm8jRskBzh9bC4Cj6Vxm5ZM5zEXx4zSLjkRZtvGduBaw6McjNMONnN05XQJQkxWYkZjR+dI5rXZ
L+QvPn5Gs8RhdYU96CHqctV2MKmCH3Kc8g2tXXXsv3XIj9MGgcJ2d5ZzgoTt0VNLycc5BDeHJYjl
uL5fnylRo3N+GWRdKyEBWkM4X4Ut5LwMmWxZ0/1bGnErDfAgMi54ThN8qbqxsWrb2CLy+6GT303F
h0z/z9melqlgVnRqgZ3eLqNvjnN9OeUb5IwSyapsgb/UhebKZAt/RTWz/9EFbS0pQKQ1P3UDvK/r
s6CCdv7dbpkKXwquCWbg4bIig5LD0XEmUb6wY+qmRcBFDav00285FY+J293UpZ5FanAQzr6z9h7z
0mUM8Ddy1LAoKYnDt2ZgB74pitUvwT6tif1o4nlcNUl77EliRHklyAGC9TB1/i91M1PMBJjfRHXS
yEJC6heVHWrM5i5xjrQticYs7h7ZZBumv5MGnipZBTzNigqQ4PuG3yA7pRG0vkbN5k/nn/ZTobZ8
dFb8Hv63pbnjRSINnqmHiSFf3XPQ/sIvUR0lQe00Lvi4ZmmKgaoCOqabjbhudwP/6sHc/w2W1FWZ
rZswiMQHSbmWagc9DNbmZ3Is6vJX4uETHbgNeCOU9mArSFp5SVa836XmuMP+NAz5FW0hm0YCbb/z
BhxwPmNFmHQ4pLltSF49i/QmLgTZ4C/ElMbf0LY2qx/TFLpIZ0m/KqBVCfr6jUbXKCAmU88n6OSr
anDscnLX1bA8pHYPm+HVNxgYQWnAPQTPcwIQvoeowVWsHpb9V0RedLDXq5Fsbjwprl3OFqG3XwkS
nyfcujjeEVqW4PVaxlWj50psuF4Kt4XtgLDtfoYo27I+4JIm4nYvvGDEmhZkAToGEdtY6XK3hPkp
yO8zLG4PooISbdduhoq/6lngps9C38O6aOGicyTRdxt+aKcpVy0jXgSFaqARrXrgi6Ci8PbmFMnh
7BumAPpZt3kqxsUddYTmwfANAOF8qQIFCzGEBEn5H6umGmj0wYBzzJxCDHRHRAVJOmzmtZAlujed
1+nYSl7IObZASy+GSZRX5MlApNS23egEQrNvugRqoRfjwfIP5X5ZtHB93CfoA7mrYRE84fTiETGP
5Ogs1tHBVJcK0U1XnK3H4gXsib8QFWf35LiCNO8EVFdgJLNu2+olIfuWF67u2DlvBEBPFxxCx7aF
JwnD11jUv9aga6uJwuNsizKZiZ9yqWsWySmb4JvW39Eh4r5sgYmQOrFeKXFDHFXIL0VqKmNXi5vm
nQSgFPDxr/Esto5JNM0L1aO4kyB8m4l8IP01/scMHn8fsGmJivhW8IrGlMgYnuPBM/UFQGVMyLlF
B0zUnPIfYR04NXwnyhn/LjKZvUZ5SE7e5PaSyY/XSvXVE4JwULOBGMTPGBJmkfCPfSPJGEAYM0x5
2wL01E4cFQXNQDknrviCqSZGifWTErxuL1/rXy3tlmPdx2Rgie0w6dFpQSZXcmvPd7zsdwwqT+Lo
KzNtYQJ+JQ96xE4NkkzQfdVPpfcTwq7aoJJprQQ3iTyYBaFMmVLjujLizicqIkrN5bT4gcWcna3X
DLD5r5ghi62K4O4E7FCwYBcuaF+yZnOJlnOMkRjjYMzQ8TFAKTrjBuP8d1nGbjpRb6iq+PecZD+H
+7zBcRDlByXGTH3IBp0zbRKARn8pMWlOH+jcXFu0LdKFPfhq1cmN587wk9W+4Y11C6wVuSaQYaXP
z0iH3uAUjiXLq+RfGLirjdA8wvI/MQ7T5wf6zGkeC1yx7zv8cyGBWED5zhqgaseZEn5i1qBb1vBQ
rc87u7oJ3opaVoqfFqjgFT5gPQMhrY7XsAvxkwqUAXzHJrqfz7HUKqSKii8rh3NPn0Zmlw9W0VjP
HAQhIxvhlKkHdRA0bjL9x5cGAR6ATErW2OH2ZiYaxBSNU7xgfN201XyfMPlkWm5f3eCQ/0En/iLp
89KJ0DpLghhRgzX2MtKp183PkitgXkYUBJTx+7TkXxcM2kfo4RxOOxvmkC+D6lGsipCZV8x5LyFY
HwE3uEoqsi29k5ArasgflOMZYk5/exVAYVkg1mb88wy51dHqAR5ddUivd4ayQJKhCjCW6vdXVzI8
9jQaU0/n0tPreHL2oiiwYmR1WUohIjaqIvdPVchlev7BClgq7s/HTYcW80Zk6xE4FiL3Uh4z3cQi
ngOAF05Naqv5Rw6QfeScny+GLkRqWT1fGlDdALCwrrKPfTIPqOzrzOTl1QQvU6JSkt7NFlflfhna
BI14U4vpaDCu/7fPGVD4pAXudELIcN29dJbLqlfQBLK5uZIZ16gTSumDKVUxDlXCOcB6zdlns14W
gWc04UghzMa0lOgn7a6psnrAlqPl5p074Cn6MxbgNqkYPMzQNwSHVzatybgLJcuIHeEBoGE/4+Cy
9ENIUJjBjM+/w+/mrKk++9l+nwy18Lx5MGYXdXehCqJtXOC9qTxP7Yp2FscmLtDYtg6pHmhvShPh
4CwuoxtXzwM2ziTvVJEMb3elfvU2h/4z2S2AdSRaOxXXlIBcgkuG3dAQkcTBgNFfm2zQhEr8P6yZ
CqsSIw==
`protect end_protected
