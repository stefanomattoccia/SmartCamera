`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
A13f8tlz6UJG9JfCNcYl8NLUw8Tlctm35dCRvt/KCTpBFIuXlOawHL7sTHowWNnYPdFQNufThU2P
nq6r7CYRfg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oJAsCu5zl/OMFEQsA8TK81YQdELnJEDcFa6KQ0EHWxmJrxei82pUrFKy5/0YZah/J8433WTkuMYX
n4DxKRAShIrdY1X7G4VuvTy06p94vL5LjcHyEy4fxae5eyT8gPJ2ix4XQa8NTiv0ndfGQZyw3Nh2
G2fKlAI5x3f8zwZZQY8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wvBGFVtHjRF0sOMF1pCWFAGskoPwO7T2ijyj/eL3cj3Mn4RaSun2E2ii2aHguV5ZVFP65oRsiH5d
RuZPDUKAsxBDhHSsGkFSPIwX9KivlJTo2FZHlBDTlkfDQbn+a3fWxc1HcR9KUBo8QndFpzMmqgOV
oDGrjFRMryCx3hlDJdU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UMkVtIsRH0SCXq8LQlXc2SFapNVFtJ6lm3Wp55oPh2JHEa2eDcLuSNAMzka2zwzCEXltR/XJthW1
e74yTmf22SChtep5vBZ+ajUd7h2t8MuWnhQAMciHkyF4IkU7ju3JOoQFlih3FqDO3aUJPcamhd7Q
ccMUMAhIvZFp44NdLzl8HbXnE1qh9bi1m8qU8jMCKESUZ7pg4lNlsQjd+Goa1H9iXaLEv3OfHZuq
AS/RQip05I1DUFL5hACAmmneYHUVM5S4EEaO3aHf1jZ3r/piru3ZRDHXxDir2Y9zXiL2oDUfsV5l
w+Pp691O/rBEAjBLQdevDcp/mZn7axrfo7gedQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BizuB2M20zTA5t6lHKGfnJrucOUdZ0HEVkxiYzkxLH0WP9VZIREBo09OejVavblw0lBdoToGD/Dx
ZN2JWgxB3v9b0Oe7EvwN3oB8w0TKm0RoqDmuPV8JuY7RwxtxkHcrVvcjXuOt8j2BPe5Ix86NYRxZ
8RqRFVGNyOVCKZuaFMVHI+ktnNU/xi6ZGsd+L0PEmNWeJ+y+7ubRYuJBTcZK6n0e0Rv144/nsqdy
X+40+rhcynqZUh14Jaqxwmyc8eu2wmo21it2TUiXXzLiWf9C/rPTasxTNu6GgF2yKIv/qtG5zsH5
iEI5vhFnzG+RShh+IHFb+FdSgnifLxcvxMZyfQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WBEZpdyDr9NfPjFUCp37UUdIujNIa897wZZ58/x9eMPhksqlKdy3SYhoDdl4U5n1JXPWIonhbpyY
qfWTq0gV9NaH1PiTuV9w+nrQziNvPhnHnWOzNrltlMQ+uTbMRquXZffmAQGphp7ekw56wGNMIqvn
BRmPzqHv8wZfX/RCaFbjfXAJEmAF89kl5TL3IWnE72Kb9o1cSvFtKTxyRoh9m9E0ghJdkhnRh4Pm
wU/+pIGwon3nUS1E00edVC7apMYbKm+8akp/2UT8ovmuCYJtcE90yRZZaeiFNpLq2UTmaGHp3XHC
2ziTOAA9fjUjv2jhCi5RMA2D0eDmOlHleltm9Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 288720)
`protect data_block
MlecvaOA8qYc6lt+j4Aa8WyndbxCWhN4VY3b3kjX0bGoZZPusoj6WzcCJVU8awr5OyaRFCeTj4ds
qy+BoWzfWk0Ws9VmBK2J6lN/GVnaWkv3ltnDe3k+yEpdTWCYTF9UPYlGeiu7TDoNptNdG8WkVYSz
7HzprJ3svHpYMOAYqkXzycGxCSdc8x7pwv7i4DdsIYNYJcits1ke6Ezu2IMUUeWEEuniZe9vH1lL
Sg2JLKMvMqlYqVSQ2ftiJRqJa4CmFp+lpBMuRRm9D7Jn7UFO3J8pVdeuz4tB0XuBPHNjOM2Ld7ZZ
yFVvUgIYFKQdkMyrIbYoMiCCGNq4pzUUTsICEi/KEm6HtzAS3wGg37DV1XOMXfRc7f9IKqy4h6pj
/JjEfHVHml3YIm9wn5NzxrcI+ax/8loTt/Rn7z5flioq3KGRVqJ+4n/MyEwWVtst1M/7NSFvCmG/
AuiJkLzHNtLXen4o9oOD0uiH+TpQswZbTH6PligIgK24kpjbEPNwh1HlfFZDAxbZahoKNe8W/vkX
TcxPL46Qh+v8UGczatlyzJwcqokfM6lsD8jBKWgANcNhbuYU7xDHS1EePNkRDScVGpWPtqsjLnbW
Po3nHvhYPbU4estahzUH/DFHN53kOaQNuOXZD7X3oiN5mH1o3K6crKfMTf7+VD9BFTG9Kh4Tq+b6
/MUJOrGLz1yYbSlK45ZkgBrOTyY5hO9grskmWTPOr2m5DJ+h7GxtEi6i2muKujhiE1yjIgtiijuL
vBKsPjJM8jYX8kVqt+iieqrqurNfUEqQcoytg+6JbhBkQjeb8ZO0mzfcaliZ+NQ6vVkfKd/6Ycrf
NqyhGzhZmQ5UlpMvYOuCvS/HpWBl1dlsVoFN6xvkTUS+FcKkWBw3+w7golzHxoreWMEFJ+ycNTQW
+KqzQP0mKyEaUjgy/Xz4YId+SnF1NHykIs3q4+Yb9pi0VRuFlkwCjpnf8p1cFolHedgtoeWxGcb7
49vaU1A6i1ySr8awUtlXW1myF5LDdZPCcz/rDhIvVIuJlnnDOJe38xI4jbhyvoH9r/QWDwJDqr8Z
MV0rky8cYMcyjsRV1SLXauy9rSPW4dKeThzIXlwt+J9HxUD1rReI+5XnbvHt+O+rL5+Spv9X+z4c
W2+th2pf/8hP+9CFdbSXYoP8EtqIM8BRhWuRqSmPIk3+OSfaDul488hLmxfJh1Fp6HpnRIGJCtFU
GQ7916fBw6+Tdl2+M/cxCnp2QHvDAPNouQW6p7VxH5tyZzd6IiC7MdShdfMoyzPLxzTtap+/EYEh
zvHZpCacQ2O3/3VLoV9ovBxA8JMTc1WqiL57do+Wq6SXe7IiV0K376l3eybTentv5y8mj2RUL0AE
nx504tpAaplHnGoSKeRkW6D7ET4aNGGBkRSz86oTAnDKZS+zkwSBin1sXEKfyJnuk74TGdPCO5dG
YRORA53irSSlecZ8LdbMAMrJWBcf74OxhKp0BY2DBX/0JD11attY7mZmicVnIlBMmyvWafN4QBF1
MTPq0L/Ega1pfGok/JfUjOfFJSB8wW6xS0xAaKfpCrzFXUjEa31tH3fMyUfueVEjEZDcSE6vkOcf
yDirL9/kGRwizFcWiBq4ajUXsMoMMPk1Bfi6MmsBqcR5b1Nv+renYnv100joNR8cI8kmSQNH/PDd
JIUlatNpsukb7rk0ARGQkxToacQiu5p/okd/scIjcLP1Pcw+MS3FQkw3M2MGMy6gPeYlSy/SAfup
NPMOCRRtIGPYDIy8I743QyPTNonv70Po1F8JECZy72+uZRjZvjbRlZ6gLf2FViJXFQ1tS3cl7h9M
nbapcmmgCVM77r9F3ZpBqO59TnBpA1c3yWx7qovqclSLk3c+YOxBGEs8itAnX8R7BZB+pCOPpPpo
5wVjDcfC2jUkbdvcHS5+AjXCJF6XjEi4uGUjxQ81963DKMajYWPccMxBO4f5DNLvCdrASzvtWtrV
GKxirlu92J2KfpYzhgYYSRQ/KBWMZU1p0ohQSBQbFOJUR6tviwTgcQCH26PHT44v1NxPSirZOalK
FEKpv3CcLRgfEprzMQMPCZpZDc8BjRAjZrGkH0Je/gdkStFvpm5R3g0uTVi9sYqXhXDvU+W+T0p9
d6J+JSyIirlQzESXbCZgETuRfnPrQXIeTKDBNnBBsyJx59RyCJ8sl/UL+8ACbbhy92sofvzTFLNz
EXd5l0RDjHRg8pENws2w8Z0mQxPH4hK1F7Fn5oeVo57iiaRlDRk+8DdcaRuByvS4cOiU9AS0v4qs
iSi90hOo6cIZGo3q3sXGR7KY/8dkS/IznKB0XL0dt+IaJwfqCsKsmcdrhJoV3105ONtZK/lyDnWe
bAFW4yWJ5KuDBSeQQHENwEQE5VrwWOW9qDFTrLBDGZdrJvcNEWzlKIsJ6fg+vMCo7nCtHDVzkNO8
fpNyqfBf1CDC1113ONmy1yioe9Xr5sgp47CQ1pBfi3QRtZJYAPFzjlDwwNYbRql+E8JIGnfw9txE
9mmajFRcdyS//f+CpJEIo9Fy+eA8JKKnBLyEuaKszTPgcYcYEhgRu6BfacKPrIMWtmpldFGWsgA8
sIOVBvt+BDNBUGQFKDOKMxY2cZo4UO+5VqWk60h2LZaDcOkm53cy/NkqBekDFrU+TV+zew/7lx+Y
AYUHwOUv+PDomueq6Ry4a2CSP/Iq5FfB9sy+ObU4sYrvsUCOjmOwbOLPn8+Apakp04IE9Vls6VgU
VEINPX/LJEMDecMp771G2kBXcRx7U6LufS4HLJK+5n24pp6u+1+OI/Nfi0Z5KVByezivlQL809zx
cuhmEpKDfASNEmIFrI6PRT4ynI4mWD/cAxgAudbGch9JOpisGm3x/fVIFPRV3avZZDqxifUkepWJ
6SCchXsyoA0b4mXpoeMv+MqVpFMFQOgkPCqfJbbGhrPHgO58V6lq516HseleBtqqEtGHL1sCgBAi
fK08bKT2ELMsE4ThqBjy13yZibEGmhItwcAC18wjjUiba4b6I/EG695IzI1rtj8IXTOqRTIebHoH
22su2aUUg9PN2IOFkhQsC+V+JJSNUjmz5eoMDKZrSQvbKC3tkm/u5bUr9v6TpxHe9X/i4ZDnyDwd
nt1sHI/70GKSQxv+GaeQI921nYkDsJJJ2hhvOCUafMQi3hbAMH8q9rRQ0/MKr8Wa1m98HnK1PRk9
KjT6PVH3IGk5P9WzHfVNNEzy3h7B9TZB99+hRwhECmr6yH5u6NKDjR5CC7u98g90w6AnvI9xw7Z3
11arPp/nExhJTV+OaQ6CiEtCkz1i08UwFuZ/1FdCGRkarwsaTAf7K8ZCvOk0JhkvpgEF4kt/RHKF
5gJx+ONtU1lUkTylizaQq5J7fUo86PjEedjocdUwrdFQPcoKmYgiMVrkEZ7pUdcbQshwhnsDMeyk
W5FDxqLuvIfnrqt3G7i7iDeaxRUpwxVUyBx/Kca9Iaswn70h2J49MHbAgq7d9FEIZMzmy7PYxOjM
ORgbYsKL+NsQlQYcRtaVGgQSaU1DAO7K/DHz0B6AqhMAUfZn6xrnBW5xoW0yoa8CnQ4agB6ThsQI
B8fgrmHeedz1WhD4aJI7vXZcgx3DHTPwVItyHAVLojv4bCp7ADjzkO2NQh2mgOXqX2C5NXKIQwOU
EVuKEpupDauM2zLaxOmhIPp+DrlPTZiVUHFyaHc9nDLvTaheaZuYyWBCUlEqmbfVme5v6mZ7v4Ej
ya97FzUdMaj/PWUQkvvH0LVz04yKqeGRkhzo35hWwESm1K2XH+ThmKBEQwS3bsVpQnbY8CaTh7bH
8sQVfvHMMi9whriDGxW0Uh+AYH8+YyxGT7q6jYcOQml3dBhlWlpEXPTSuwZQepZcj6Vrp8TgNxX7
OXQ2u3Bh/zYOE/wwYn59F7IXhtrLi+X771DRe9dnREdSI2KwEKMj2c64x9xG65iijADDb3A3B9rm
ntwudFmT/WbP/wknYZaaT7tfe/VBrwwoRyoPDvLe4LxX2On3/Ywk+DyOn9q7U/ATpN8RYOSX68iR
5RmHfojngJPwvfMjhamNldhyBiMSrsB9Um3CWdeCQgA89GFrm05Mp2LAynV/0te4gG5UQklSUbPN
/6v6p4+jpFmNpnoriS/kJ/UBTUaQ4OQV5OEpml3VQ1tysHN0K4o88fkmDRW+582ttnFWnEBj4CoV
/t+IYAW526EP8DVHNxS899nO8lVlLoPai2bTsANkGs2by/Fe9FSOCWIj6jsmCpLyF3dxgibvW57m
Xi+Rm6PWesLMLxpM3y28reWR42SNXDdBorpkUYUxpDF1y0c0aH8z6nfl/4taLgTdxTaWDG4weTx1
vNN7kxH/MntVgCpTa0jfNneW5O9xfdE1kFLJ+Cu9kTEjcWwNwQIwyiv+RnKzFW17GmY2RpvLt1kG
PSV1Ld3rClrF8tOIk6CQp0AfaO2eGKbKVv9MiPA+F0LUe8yJU72+eU6uVS0hi08Dco0du3NjEW5F
oMT83VnuQ63jsSwAg8BqNsFUjVOBiApFsjWorBpf5F55syUICCpbVO5SU8/oEmH3lLelptzR43EO
1qTUaOZk6w4JBUP0rai0M+QDDrcOTqQ3dogW3Y6KlYWp/Py1UhXc7gPIJeJ3oMcTv8NnelOutZxT
cYwxkdqVtbW1V5M6ly3Rw04gL0P23WbLDGgZ0mrR1Dy8CcnoN9x+OMPa0okfJDPYedXoYw0BV8Nl
JUI4JxJZWO1hANmli3s+8bBGUVF09XRUm3gXGiyspPXBNovwPd/4qTqkxyu9R8Ht4kS9C4c5OfN5
DJcwGHoegfuUEzDObV7WgluCt0eRJ49OD1AND+CrLNbmz6OKciB8ac25c47yxTiMrhHQIgfCJl03
cPPji8LPniqk+4daY697Xnrr+IMJwYJ/X/SgqK1bNFQt5NBD/8oJ6KKgUKf2lW5RkgHMbtz73e2J
4csNlJwBBr55F31i/B8aHyzVw0/kFy/feEfK0I7/Ic08IsUqfC+Rv0ZZWWyf411z/1mp/AwKsp1u
vyZIrtxfv4wcAOY9EtlzE4SuZ42nKZEFjchaRs/5OkwZvZiR0w/cqR34RDs++Iu5ykH9NbEozfoI
q+B82qImTm0IbK/ltTRUvXMtReIUk8UEC6/tWqA7toi6ZWqa/+1/+EFHjtUePCr228YW3HRCtzDT
nxVYRfcc7i9uKhdmoB2BpM6HZpNY2Q4BZGo8wFGwVQXENgkH/FOGm7bSSjgs2FGqzcgc1TWPpV/5
vZRBZkLK43Om8OA1fiFvyeR+qjSZF/TOXuSVil7emD9N6ZEFyAp1NfSXlAh+0We9Aa7/VBRRkLz4
j/57KfdoHthrGl3rwK++zeNyBNb705/L9yGZ8rMxr8+XlpqXcUvo2Z71Z4X2lSrWSUx5lCIqU07G
u3ZUycavVi/ZR+d6Lu3xbirk+vr4Q4G8uWZ82ZdiKq3b3AnB9TaliCtfRBeXAQMsNvgV9mmWFYja
3pA2O/jHUO4rJaPn/lmqic8XpkV8oMexsuN+3Phn9HvYK4TM8fJnY6sIDsgcDILQvrrzTE4aAh8C
QE5lojiFjT5rhtpv2zXCGUHbj0ItAs4qyyzh5zd4G18rQ0DXFO0wb3q5cSekHjewMdt+TBRcRPrn
uLV3HKbW+v5u27KWqT7FWR+4bzTcjHDP2L6nmVR7zcdao9GfNjVrzBUXUBgx0nQ8q1RMkIyA4wXn
wIRY6M7MXtIwhmX/igy4/0HwO1ZNHlZwbQifbK3/nFfT4wgmXGz6nQxsLeb6TYpgYgUwbKiIZQhT
tO5KvwwsLsRUcFgsXOytaTeBgW+w1T1dn+gYrSzuY5exoGtz5FHdS48GxW1XMgiw5jydXb5kGL8F
J6ftqlYOrXhYboXOrXVQaOq5k7jYYZ3Y5g+ry8iZhylsuuseVYrs0fZtoUKDWNkExGLmr9XgdhoA
UXBMU29J9MzrJBF1TirtqIptZLeamgSrsZsv2/oH6xKqo2jSNzeeaQ3f7QnfKwJEmkp8kdm1Cneh
9PvnewH/QwGqsG3ubYJ1KT26S92EtnB6CI+7g9Zvv3aigqv2gtuqvxFjnhqgwdRQxHdXoP6Bw+O7
R6Hj5rstcyx/2qDMlCkp/IUEEkaAoO/3JCwW83QkcteFgsDMtqs5zdtyw1fWHcqmjjkmmHkhYadn
S3ULCkXPXDNTG4fzN3fzF0ojSSgqi5gL16lcvYjgqxfwYzLaXdgXCc1qfwi/FGxwIxS6kNgjGLVw
IGupQZ6caVdypmTT/9cKbQ03OOFORcerQgH+EL2a25kzudZg1Toc+eYWDzg/DypWBnjl3WQ+HIzL
HuAb23wKZfqYPHLKMU/kL5nwIrVbusvH/0T/HXjHTAbKbm6lF6unKkbhubXJ8i881T8QA44P4iDr
hB/6PYFfbp4RSnjiL9Mlxg3Zaw15U8EjtWnwkm8rQn9bI3YRLPsV+B9bWNcr688HPyzWQMoC411/
QQbk51+wkMu4i3+jeartTfl79OQgxD4Ua1NWuexLF6pQ9BqhFw6TuBpsGbLikef3TNUScHttC+Lp
iCam+pLWrevWHERPmpJ/HoCuq2a1XfLCDVdv1hfyHmW+Zq4miR4fx736nvYDVobay1Rz5oR3Vuwc
RAQluKrVHqeGUDy0CAN7ws98sbh+1A7agbkpDuHn3F6mC+F7vexZR5cKGfWU8N+aOdlydoCU6Isp
sZBwO7vVRtePpTOefDs/Qum8FS8m88R3CT9ieFdhSolOzZN5NFujXJFuXNaXElTb4HCSlQC3P43O
8f4Lyxsj7xfUez3rl44g4oDauynY7QTDY2ucjjaNn333WhzhArRssK8dxv8ggjtrgdCueIie4zES
Z/3B3xur28UnrM3HmjXv/SkaA15u/irOozSLAdI8nbeHuRPV2iPJMt9u75dbAKIssM3ZYnvW3uu0
WPF6iwLOrCmjOsy3UROsquhDaqgXNhc6DG3z0PNXV0rgzpvHWx89OjxhrWulSJqYFuQFjTp7BLMl
t98hLZAJ6q7pZ4z7g+NAsyfdwtQ6DT1vOcVHfdTFo/JpGauOT0p7KH00b6rr4kryg6kcJe9c8zCs
95Eo9ZdgkEfzshzezJb1s+R4eh+CvpDY2dAj2mI9c+KRXKltQhxcVuGfM3TZDPVxt3YlUD4d6hf0
GRYTk2FAvNNq3hkEMN5HP94sLUn1+z2wRhfpT4t2uhQPJkMgwK7WY4Rslbrywg27Dt67JD2/Kwqf
Q57Y4UUUQTL005V4WkRdnEF18BKPyDV7ksGBtrLaoyzdeA6xiNvOCMcaiGxzWo6bWQ8dWOY+CHeW
Fgq8duw+kw/6BC8lSS6kmgMuil0SPGgId/cnb9EW+gS/8vbiTpnnY6kyXjYsySupFm9V+X8D0rqp
NxvtvwKI3WgTw8sOd0oPN+2VAtAGY2Lp7ZZW9DbFJ45myPZ22wDLh2oYalHgLXWr5Vw37YZe6tiz
stq2hrTI26mQfJXQopvQRoGGF6QoPhDMEFiS4oKbb92+MrfD9z7Tgv3vpUPpojR4/KUmALxv50VA
gKHTW3JbH9jQJk566nuaFX9KlZA+eXBAfFq9sF8a9Iq+zwXFBAYs1EoMNBg4DIZ3U+nnxpIGOpkr
sKkcjSC/ZqKkYh47dggIqQnTB1ckkOGuYM0gTgJSdSxd2Vr+59oDv7FWXGNDLP7R7kjdlObOWy1a
kzzYOFMJqMsux2Oz4v80FZqtfFhcL4F4Mix4rEhvFSk9rZDWj4EA3EoC22/iccz0LQ1eZjKlLTSB
vekzPkpcgXbmT7Ldd+Y+Cva3TOiU35I/C75e/uvMFfU+Bxuj3b9BymAqZNdbbfq97DCI3kdV2813
f5BEgbdSOskIdfrO20+jH2l3SjSj/ZSJd6jCIkx9p0KptFW5XSNumN1d0X2/YOwYHQEXeMpSVzPO
KFAONyO+IJ0rrmepBinYbFCc85dcxt8PD40tD6rXu1k0jH6uoJX4KQirAlFGClgRSfEDNOjstHbG
f0abXIISndnZjgHlPVw3yHt2gjdUMM6JSF3iAYewSFV4pVwLyyuo3tXb9zHHYG7amuQ3xndBDucZ
B3e9mnXeO1GcHr+8gk4kBxtJui3dzAwrDtHeldmgl9YsAtFRtFYt/dBb7fSM1EyTRt20UXzVY5sh
y9pDp2MIsRjtUc3XfPkLGcGCRBOsTX5m77o34KKIhP23DCgt2sZUK1KsOwOhyKC+BlILCQZ3Tl2x
37bZlre8+nnHYCok6k7eM2jKETIzx7JDmOSiep8xMp8dw7X31mVgSYLcgrESo/4mR3PypiPqSkKO
Jm50xWA+t3widKOhK/ovEF7NlBSQaVBwozEB+gd39wD4idExhOEvaDjQe21wmbkyNSIu7XF4koRW
Dgb2E8K+JnUEgJTH9D1bz1+qghrnq38q2Ard4xbjOJcL6YHZyd/cBlSGrEHUemOzuHSWYeBwnkkq
VaBp2ZSF+TX+VB4i+RMuOhPnSC5HB0uxQhXcUQjS/qAsdzVFOPeccR2dDm5NGNnWhQuZhUtWfEsC
Gkqg6Isn2tSYJFcEH3CdKETM9xrQnJ2uxsYL96aYZEaXtc/KMc2asRDmQFPbxwKFn4X303r6368Z
kUr6K2hJH4qGRJmqCCHLAmH+Pan72oUvNalLfwfvI3JvV6KMLn7CIgxEx9Vw7ukzPUr4WqKptlTS
p0ldqHrDihdYUqPktUr2w1JUSn7tv7FgXUN/1AFFCTrD0drQzu0aDUbiJCxsms19pBKkRBJHkwTJ
VK348a3rBkDphuljsykBhbPMBmMOibDkPkKgZAN+5XRuoFGO2nwWG0Hhvm1q6YGy6ylkuPl7/NQw
65Mm2TD0uJqGwjZe6u/EDHTEzF5JjhZhJicdfFrWS5jc0e0Li267e4FPKBo044eiigJ6NaEcQjpK
oCc2r8OI984z92UYat2NGgNdJVs5gFtfReYtLpgbZir6Nx7RxeIBChx7FPgAJjYMGe0Bc4MrCubX
rRrT36YxDvEOcdnc0wQlCTEBOJMxCwDB2WJDnD4LxthFfwstQm9Iov2gYoAx+vKFntKaC5pUCzHs
1zPiBu7fuU6pr4a1hy4yeJ957+932Z74d9IDjeGUWxV6sstJO+eE8/ZEssCyW5VdQdNOVeFte8pQ
unF0tYtP5euz8ZpdLXxvYZFG8vUpMkjmuDBL55FBKI0EGSLji9dC1/Fa9hPDgqZShtfgglqWNu/S
+xy8UiUvLT7ekxFUCnu5/JWfhAQ2sS3PIByEn4w4wJvsFVRlMLxXHLmKtg/FqYfUlyw9C2SYMGJB
63y9mQkBVKqeX4FMAqiiKETEa0oOHOJ7pkSm3GnTJAJSxNOvfVwTUKh63C+olmNAx9sXNhPF1GMT
UPZmbs4Kk5Ow2ewTmSEhMiTMBgMnB+Sq68mUy5yiLfvQtryRFeKjGTGcfgUdjEoch6Nk5/6eocT6
AWoTMBEUP+TnZRWLCwJdws7Nv056yB0fILUlCdBxo0gKlkAPxalTOhJ4losgbt6XDynQXSH8GUqr
dmDp5WlrMakpUuvHR6c9xK6FuRcq0HuJgMDCUm7KWgMnc+YSjBzp6YEXzD5B7ikywBu+EcGjGqZz
9kctFroPDgQ8aXpvN2aIadymzKtimRXh2VYfVkyI1j0xYVWE62azg0DfzwV1bMsqLkPoCHNtKOqj
/fF/dlmhCEqgb8AIPHKrg3ImJOLjPDcptSLU6HuOFi3IbY7JpHq1s2/vNGpDdRRx9mUxXYDxcpYn
kyW7LcUA9DJCFEILVTP3CC76c0js4zaJ+uzfND1fV2PsRpienkQCml6l+8OqSE0tRHkpqc+owx67
Hf7uXYN985TrEHftpu6HLMtehSA4EZQ04v/pUnqyVUMKsRfvRbFMRLKNd+rp9EIeswQJmDrE5WB6
9C+5dpYKbrBDgOGJIHbHO8mm5BRmbaMCAb5oC7FTi/O1f8xl9/XSmF5u7Og/GzVA0e9vTrauxpOP
zlqdK2nb1UkzJI/AEBH9wcE2dkL+WuGMvJacS9I3+SwN7ki//Pbh/q722oVO4AosmxpSxc44iLfR
TQpaXIRg9sXuWOk4DweumjSWuUkqJjrkuz1ovaV84y8i9T/+4wLBlBhHHIWL0GJI2+6cCEWkpm0t
m7wwBEMVnJxd3V/SqQw8qtcVwPqg0kAR45geZMM64iKLjQh1Uvxl9cPMbqF/cKYXXu3+Erx/pf/I
r6SSumqt+cqH9z3Gg5+MHEypiNvqcKXyM/4ogbFk2QpdoOS7Y6enBUsFrZsV/YfrB3GzI/Bt7//E
Ie+xpg6hhc8JN6CnMeemvlo/xTrynbfpn5cLK2au8e6M3mnmserTRDtx1SPPbU8BQC3uzLARYv6W
/fkgGu0aFqbB2SW8UYSfwHB6/kCXg7sbMHhSJbzkSV3KlF4Q4oC2d6BCgg78PNsty0JoAq2QuXhr
/9gV5t7aHPnNhlz2c6+wMcoeBwcbAqXsMoL63CUqiXde6ba3uJdIXfRBlAfthenPUNtQve9vVJlE
bxDBhPIz1dEg0UWmMenBmbvMaaEMNkv1Bac6LghTB3A91Y29kyRoeiWz6roarH/QFFM5br7DewB5
tY0lKZl0ciAZK25gxZRNCsWBJXNQRos3l4J3v4Vns1zLvyPRUPEVYE+0Pm/8ZRwKexE7DMkSmqN+
K/jgdEXXncHirFzOCcOSDxuMewqolf+MPTxIyYR3m1CknPMVCnqi7NzAXzQuDFO1sDlvt7RbxFUB
nFDa9QBKfrC2RzdGJsDZmK+vGwiP8lg2pcfTFnzwnmCOM4zwLv/WToKCOj7vDp0zBBoH8/Slnr8f
zA4Aq5C0i6dbX1K7k8n1jsuF8rG1RUcrWrMoSh1jM1wUAoenfWj1p/sWtdTk67V7d7+nNEuTYBMd
/oMRsF1NSIlvKSX/8wkiQOSpj++DcDmG+YWEOyoe44EHh+wKHm6sat5j0LLV8uQeaNlvkxQl2GYs
mF+F0W4NvxmawnqrHvDTR7GDKgmm8WB2UHgFCi7TrMe96rG2sOmikNrNL0b7H2JP+Lqrgt3D2egU
kMy3hymX8egu10gb5cYZaqNoI7fZDCv3fD7x1MtNZjg9c7vDYb4EzTTDfTCdUsxZjlIEv1j8l02C
zmRwzkPz5VhGh18f2WAIEm1fP94DTsYQ2So01UqX0Z6hO9c8dsGzgmHoumCcjJEakS+25rrcz3Qr
g8JQvSiL0vNEUuTZU2TIo2bqD8ECqKn6QxwsqwZZ9n1pNwsqJo8+OoRIstbc2mNw7dbo92+28AxW
oUOq88sOY+02DlF5pVO1/5HAxaDearfo/cZ0adS/I+9YA27vOfeYp4ORIlF/VqntXaeinrKlwO0J
KZNGhm20o3z6alcv6Hx9E6AP2PijB7HY7O3AQ5QfWuTg/XCQFk6vWQV3Z15saDeXZz57i0CTVSIu
xAlyxUIaWo3uJ+AUoMEb/VXPvLbFEhc61x/ZX52uUVV8KU4fq9IkmV4Qxywigl95T5BtWPYpR19w
4RURC9AfonDsvaShBnYXQb04tXQVavY4MsAPdKvk2yu2vCFMH18+pG4YlapBV+xgJBh3SfOMd7P7
zFPjbIBI0MK7jqktGCQ0IgV+2wpcYsuODj9vcMVjITPX83xkM6rqHvPsoKXV0ApsbpRuxXrrYwh8
GiXc9SG0O/yyEdu3VVImjVkXMCpJ+lEvKsNxyG5QwyQgfu7Bk2cPE4QkEABQbtrZ3EuqsTdgS4hE
O/MzjJy3z4lp9lV/CYETxz8PZEuN/0Fa1pIM3EwcPAkO5KKD7VtqnLvO+eelQR6Ig1g0zTJMgLlu
ayVbCUam3O7ONBoe8M2FRV4qaPSD3VHiQJ3DpJD30rYumktQqKLn+Im3O3T99/rWhuYMYmNdtMqs
bIJhlJk5RtqW0cGpSPDbysNtc9idu/pgrS5E0eiU1Vvvt4k4s/C85iAwiPEvA1Gfx7lWKrCrvOsr
ubTczIglBBnh3ykSdKMFyldECNYZ9OzxNVGhklICTYIOFKZmRUPbB+7EOvJo4bEEMMMMREQS25nL
f+SbsObqbMrJmXvKkIUaJf01M8gZNEZBP9pSEGd5wu4B3b7jLC/XUUPVuq8j+zN6CHMaVCh2iQ37
RQgHNqlyulHOPB8iEyhvQ7zvCLaWgUW93dMQqsxkNXJr0F296sTGroTulwg4JR5YiSQp3y1JJK7K
bGjcqaJjAmYp/hak7CEOaMMTknyU/unbp5yYSzn/STc9HihiwtURUcpWix1MJEAZBIrNCBNWCpgM
2jXhrFq5Snva5H3ECOou5yKx1pZjT1ghZiXAWk3cbNvwQ5ekbP8OQGU6VA5hdkhNXZGEmV0IzmVB
PA2mRAwLFCC6gv8bAR9lY/yTPxiOvivvB8l5ATq3kN+igD1J3XtanjLbidIjkv2K2AdloGZ4pqH3
LO5j/jEvpQMQh3QMev40y9fMoGRJtR/oK8djxTO4m+3hQHPWhaA6B0xy3lQM4A8l3oemSE3mj3XM
0FnhP/9hObbYjMQwonGBi5u7lY5ABDXx6Y85ZfDEHmj8FtAVwBStaa8+mfG2P/93Y3Ptvt8ub7DI
enYiVA8dlY3Js+g33F7ajF0/mRcOvt65h/l6bSLM12kTV96yHKPV8eXuIuFejIg21S9y3dv1ih3L
5a811ejXPROF2D2uXnDsMyou5u2/A34pSAa/6XNDQygGRgCg1nwvwWMOLoX2vguAxt5SbZ641/PV
zGGXAt1NriNxcndG/fMBxavef66pVa+Nqrdrerd0BNTsqzE3WHNIRsAe5L6qFTP1ccwRX8XG0EI9
XGcYikdnaFuw9rsJmCws7Mu/B69pj1qrHz0h2zX2k+s+B4XYkb5IbHpSIMLC3/IQ1WODAhdoqXoj
jKIsn5RPlyeG7weyDdBF3FFgzHA+z5NSiVFXP8X2zHcUz/0PM8kNcSFNUIq+9iUwxBL6jxvtCleu
3os7vexnWjzV7/hazQ2wrqrjebJe9tM8P1gJ14dVrI8KxWaNfqkjSlUBxpwF3XtUjqLQ+QdOwePt
9k/SaT4l6hWuoG7ZeJQgiJ3toHqYXpYOJAvq8uCQMt4NQcH7rDQUFte+nES+wZt1vU17yeoqJCoi
JZc5JnivB0IlIQGbCqiY0frII/2nZLeywW0htn+WhYb2GyIdwmIMZE1/r05vSqbj3BQX5zxyeGld
Ht2N1zBzP5AX0ZF3SSFlO6UZRy/5QoeCGN9ODBXRm1a/qbtR7eTZuPJ/gab7oBtiNjg2NXCt7Ol/
l5u3ZXEhqdWGD9vZHjtwLw7YIy/viOyFKt/X/IK9PKEgSrXwxmA8AQ+XP3EiH76Lnt3BMnFz4g1P
AdqWiOA9c2OQ9u5XZhckbVNBTk3CbauUllDYoCmfNMheOVEZohmOGo5mTye0z0Bn5MRAFyW3YbFn
qavtTGndY+VcjWFK5FbdYOFrpZmUzs2TmcvpLftjGKxqMkP+f4W9RWrAmNAJGR3DI8mZXHWAJBsr
X/kwTqwmAscW3cyY0ARndAVV3vI9bn8fV7KY13xNSqWO1V33KL2iFREjcNDjhQt+YMAxjOhe/nBS
GZ5LCoFQwbqnIjj420UY0acXLTKEwlrKvzqlR5nor3tfNK8U8h6z5L58hz9ybqMwUdJpYz+F4+pA
Z83OhpUIstCK3w2cOvSOwBye1R3vlp6AJVpE+e6kRMmMSrAFG+VcQIWKiix0I1rgrbiQ9IMARcrn
0kdRcRFD18nAQge27OFmwSmDuXhVeylhg1SBeJz0qgPgdp5A2uFAb7TLUCLdBejLbKgf6RSTbg+S
JyPDWf3J0dww4vAXlK1JF/Fy4eNmidzolFBmIKeDPbgQB52lipZGdRo2oXBMSTlAn7CjS4/x6QKj
6kgwDdlz2cTPE7ZVp4ofxhKm/hdldVZtmwGXrPtLhVdZofE+ZdtKeWkt0d0RYRoy8jih7vuPVJpZ
0cJq+PkYSPAZfTci/OauDrtwVn1aC7XWNHSELeycrYKvS/IN6Xa1rSxnkFNFLQ6dyEv2vuM3OXdp
2hvDS0mpksgATXihK3ssp9bXS+kd++VBhw/SF99ckMqBjVdxJ+OOfaBlIJpZitoBgMMplN/asln3
qYuLAMnerE09GdXAkoRWGRK/h9slsTFNrA66BLajtOaNXKPWh2ZkxruZyXzmjv7lssK62PWab/bf
Rl+UAtS4jjbZvtV1kb+19QkbLLQKr71R/8wdJcMarYaNk3LO5jpf49hqVbCFK2N0GkkgpFhEjAUQ
LPkL4lPeZmtSsjP24ilwtg8PpGP6IVrx4SmMqfgBKFnftu41PQEpzNdwTzv1/jLp9n64B/jtS8Yv
OO59NJhV6EoUsquQuliuiHxaOUDb6IsGcAILYKtQYdd0SOcYoeLkifJt4NdbS9Z29BaW/Duva0Ue
GOF8Aet9bnSOOtXmRnAgaFkZ8WCnkPzJBaVKFV9kuGmQ3irj1a8S4wfJ3L8fFQZsLWs3HAwLcZFE
hoV+G48OsKI+oCJfpUJYEE++XTkkk1Lz+/gjbUwxu1RcSude0pocQeQ5aIiKIeIiPBGhbdSwvyaX
VgpifFsJifXuX9ZOPbTdPQzBvECKlXsHp60rpfy6i2VqON85+qsM4EWRGVSkDcyGblrHSJpPX8BQ
cHLM3Po6HeAcz/DGJesolbtvHTUz1fGFwKsIWdJDXwoisDjPXabOFxbp6Y2rMHELEPeFeEImtaRi
htgJ69NXCyy33/aO2GJKJY4wMdDo5QGf63v7hnQQuxkfyJI/v8wiu0ekiL9ZK/scans5nkEMQfb/
8cgIaIi0pB4VvpT4UidGrvZVNARlUp4mSuSRB4KnqGPUh8LJGZT+AGhhx4yM1trL8+Co8DBPV+uW
zpreEnzRBKYRpv02zjxxdP+YdTzQq9TK+uD379kWej2vaBObyr4KZEVYTvLtu2ho/K5FuaR9rJc5
EL8zwrBoVf18/JIuSPzp8y+fUGROxt1Qwz0L16+xfqQFTI4zf9DEp3PlZUaPv19utF1scRAH1W0/
bNxFfyUi4besKnp1O4RsnvSgftHuwh3UcaXd8UOaa6Yp+8hCbKqHYqBiW7ODF42WVV98ETwgH14a
IXm6hnCo2R0q6TqCqoXsg7L/4YNAYaEQEBEetht5WFsi38H7Jwabuc4RiNUjwXkluPq2mBwZbKgr
2FGA/x0EgqrxpzqVBaRjPdu6sGPSacdjLtiVHu3zIzEtfKGTkgotQJirAvAHDeNVHDnHUGhjygee
YtqpdkYOMfrCHwUleSvR5hD0W+hWbl9GDkvOhDOyactgBtUecepa673MF5Ld0HNNXbAWnvKBe2nh
d+PI1GIwkPccP1C+OybXzMq9GC3JG/qw4R7clU4vC2fhO99TcLbuVUc0vnFuabUQCMrJ0FsF+pm1
IfZoBvVYxvAq+Y41d8rPQNk7W/AresUOAwOzsK514ISKIoTjPNUs/Gmv20LFVxqAXuEcPnNoclxn
rHgqVNs+Er+dXnGWc4B7mTWeAfcgM2y5/uwaaqOdH3Z4rky34vbO2XRLiTbZKqu6w5QjlYCGnqZj
0LHoNj772JDPEQ75wWok0SQg/DtWuD5Li7bukf2GkDUe1sCZNCG6Bq+e3wqVKixzn2COy3M7xQSE
vs3+lQXx9b4kfvshryWpts/SwGxFLpIhYGXv8m6k5HeaALLQ2KGan0Pj2RYa1tLRYaYzgkjFUIFl
ZmjkBWZ63WidLoHo379sz3qhx+Ss3hTIZ4Vi77mLXu1h6xJqF5KqC99RgRe+5z215DaE2dZiAKcm
NV4Q7dxdAmqc98saU7SnFgkH6M7kTVuflLxyHDLR37hqQoewfwTyHbqQirXroggc4v77ANHAXaAU
FCe2UA+BN3D2HVcsnCQtgahZjtMpbmDtF6oOY4/bO6MsJU9+Q9A41uW3H76YAUhOQs3JlXGvGA8Y
+RTZbbhtliVyc8bfydf9i9vazEOR6QiHMhhB/ggf6rnP5eZmlvlvy1vgH5NQS8kosf8MOtMECL6B
euQPlUxZ/sxjek5E36hpu8NTznncZCmmQnuRjl4x0/Ac7VRQpnS2pZxQWxeDiMXcZKIYEQQwbF9/
ZRmIoH+QUtV6QKvqAr3Hoi/t/xHZ1M7H19iPA10uknksvg9B9rPcB85Mxjs6YGbZhYmplh1obCum
nyTT0tUgSeiDhu6aWsQrHpwMNCio8cDB7lJ8Sg1VwBNN1ISbkFDpGB1TZ8cIHbmz01wgilUGLiYe
GDqUzqCdY4XoV9cov5WJYbsC1CXCA4aShUXawGLx/Ew6KwwmoDmVMlwiCuUcSEMXxPF47JErrB3a
vl57l1N0vQCaIUmLWGvpRLO61u10b7WUsBdJuiU64Bvh6QqJ40c29YabwgxksT90WHzrXJ94802o
+7hArr/RvMDbR9f1o539sXtKGue5bU9F8DES9M6kX86DWgYYfAhdEsGlnY/gI7VFC7/cbOaCMG5D
S/s5ONt1FdyMJ1/FFfJXcDXpzXbmA1QA5tB2iAa8UB4OeV3kXZkWCe4zhTv0nDl3I7vRDbmyp16C
FMQSUNkMvEdvMBETGfTmrAM9q2d3+kBaCBz4AZ0PejdJg6ILhTwXsrn0NzPx4IoMG4ASlVXuhpwS
9fSosLJwIy0Zj7j92qgCZeZPyDHspFKYdvcrfM3fCsYVaxz+XfceQKpp86cfMLrh2gBuOcs3lBYt
B8Utun512GisMJZNBEDChszsQUBVADhOmVVky9OHCOqO1Yqe55Y8R4P/IwGLIwSLz6y6YX4FAepO
py7B4q6dUF99FpSwwwyHEeGNNkKMHNLZlqsx2psETaVCZb0bhNJORTg6NOk9vHz62Dlay2NxzHD/
7akSMzN30ZHH4tEQl5srGQpjjqVk8z46A0DrEdtUUOpKyvuE2XVurkTVb1s0JDhgebdkLsJ52Dsr
DKyHfRqZLaHmiyHNiOwQb1Pi5JLdJ8YVPLMHTtdr++/yD3sVIQ9c1trdb0t45HEkTqrokWs1YOkO
3LhGZfAcYwhx9Af3q30Mq1Dm6Thrbxwln0S1/E5xVfC+viaBDQfVDBO2+5YnPwvtedD5n7MCUH3S
l5v8nF5mbFaKj6mn/x+TNndqUGJKYECUQA1dAIMTncqaPooGN2FFN+cQeptRPrShP8xRqLj6ih8v
YDJBZkzaxzUcV7xpMSPK5f32aBQbAqJk1yt01YUJzfxx7W7u7IjUgpTlHbtkfRKeeUHicunTSEFm
b/Z8XGjC7zs5tCPZUbXeeyo61XYQV+honBqQNGxehfjmRC0C6+KoD23I0vLVAfL/oTnY+l3u50U4
Ma2Brk16RVt4/PZdW0k9AT7DP2KCd8r22uRRHPBHcevUWTGGtPZemk2fuwXAf/xEhi2OdEc9n1Hx
QCqlbv0TqFuhvH36l42a2M+CYeh8JrlW9mYaOn/LhzFvKLZRw8/tusgUubbmOn6972cHAlwKCH6F
1zNz2oVhc4N1nhBCEZ9T3p5hab8a2kn9hxe+gbRA23RA7nM37GBfj6TH2woAO/C4FcsudTs3wmyW
nJJatcL0Oqb9mihCVB8/vxrU2NYc1i6LJfAhVdpt8xj8vO1uxeLtG4jwkR/aPAO/QdTrbwaqo149
YW/p7tiIZm3B05c3k+mhc0Rs5ZMb9IAeZk5wgK4cqLrKyJ0j7YqtNZgbdjwPfxEhGZuWaY7mYR9V
FX6Y9WyEx65eJ7Kwc+jf2fQ7xTJ/Ghn9XTAL6Y+/ldnZQ+eJ8JKaWLEtG9ZjnIOzGA1N6KbCYXnv
YG7KBn2YZQfU7tTC0dkK8qHg25Gvn/zhXUa7thZzWdI8x+opbWbLYibK5nX0OabXLTBzaaEw6iS1
3/9EGi8xPMvT6xXCsTWZ9Saxl/1G7P2iVHjwI64m8PMKs/qB4axz03CiUxSBF+zj2D/v/ba+hR0E
zTUmisxncyZfAj7+Q/cTwUJEXmHB4V3pM874+qxxxcPCO8FBSfs5CuEvTp3bcbS5b9jJkEnougCZ
VJk23v7HfigCnzAwKdOKRRaSbZXJ1DZ9d5vDNYRjDpblR/Y6EiDaPQynnQOR73YLjNGKxyJpJ1S4
Pq5OGq7GwFSWuZLwndH2mG0uuvOtEgND418bL4+qM2WY7F6SQQ/DFEyaU1v/zsF+R/CkWuwbqEMT
dD6wmclxYBSzOIYBU1/Os/wuo2UWoEphcicpXp3vQ5rvZGgwjEmAQyapNm1360w71dtVDWzwOf21
YwGG5J+KbcPNQp5KCv+dT4HRbLb8VCm1N7FozA0LPGq2J7Pc3RibyMMl0sFQwCTD5erFi8xnChck
39f7YIByKg+P5g6e/ODc6wIgNdySB6sb09HhiPP/FIyoyJ2d/OcEvvmq55+6bR8YGi7SXHMCdW/z
zgv+TOi6yq8n4240dvQgVOwzpCfUDXQrxh814U9B+yDqI4DXGLFlhbp8uL/8c0KD6nXfxadn2VsX
OWnlKR02LMgeej6t35mtaTyoG7jxzbisQO8qYJ/OLBdHdgqfXJYdHJ9QDg0wzGB6Xw8OpaKqNRm4
7l+sbHPf2UXDUUeozXFlcEekX/Tr10Gq6rAizW5/ustMRpWEl9RntroUmuCnWjgbXVQ1HPJc8SAf
sMgPvBZzpWG5AUh7U5P9K3dtCTUMvYbeHBu8sjpFhk2sWf4JxjwqU474S2mRbSsZcnccGEtkVcYm
NEG8swANnO8LaGc2cdDo6LYsdB0sPk6Vefv7S4CtabpQzIq+/CyqJnxU5gvM52Z1UaZBJ5pEoe8E
9DBO5uNxekyUqWaOq+FQgxZqKXFuX7dSbHI+woq0rPbci+IPfkgenRc9srtl1PK0eUS9E1y0HRSk
yzY1/0GgxmB0Sk/ccGBPwtBPIF98XzTTlFrylqwucwrXr+bDfNdLQu2Dyr8m73TH3tLP3LQR0Y2H
V/SrnQJf6vLEsHQQ/bjrqERp0XauKOV10waA/CKbaYSXPnbNmyVCRDyPTwQnagzGnrlpH5SPgxuU
0NFzRzWNFuKXlHJjKQHf00aqmebML9mQeQ6etKVFdPoW8Hs6hqhRUgLlOejqEtFiPB0HrRl6EWKW
u6lPEfk91K+OuvaZDZqh/4Bd4gVs2yrSzNrC3E9/g5+Fh3ixSELuleSw9P3hF70yO8RywLPe+Xgx
35CWQEEQS8QPwS4wOQi3X84/KJP++9cxHFEGmbxKTb1gHcYd/vzbtDPO401YZbtt8PoFl+Idvlbc
XvVgLm6AGTWVbLi85/u443AgOM27WXmmlWIiGiKJ3C4EGYg+sn/w/3dHK0EjKxxTHoDDwVy7Niaj
KldA16B3WG0IJvOIRxImeoUvASQbTsDQyeEtl5zqGsBaGSNTVsR9qwgAoyOzdY0DYnrhwjjdGKkE
XHXtJ/6odBQrmmjaZq30B8MxCkTjP8NK2LWjQmqK5zS73Cr72E4fki4Qmym7GAjpsDaHHlMAekBb
OQhokzwKIpE/C3/qHTBBtKqFXBu4hPp45fyOE5h1jGA/p9KJuGizp5PNwfoXM/Gu6KSutX2PQlJa
4nVAtHPFQhJKBg0NvMoN9wnYRFKn29CNsCOAp+U3yzC72c1EdFph/ww4wdMSyCpsT5ygVsZSSfRi
ESL9TLv2rxutMWxeqJpD0Sdnhht3WgKXrcSCzS7FYMHtK5ZmcgW4TyfTkyHkCkYUUoD/ckExCLWu
6w1XizQkFbrHG7D+udk/3YhtAcrNYfJPt1lGftI6OzNm52Ww+VD7Eemc9WyJBpp4DfQlFX2AOGxf
4QjPbdgMSi+2oWAkETU/dp2nxwQmCOoFyyoK1GBM9ya/yqPkJzn6lH52utPDS4kHIenC0oxmNNad
s6uX4TUgmXKIMgy+hkeTzYQtLoKdOUK/iDQn6TlB4/JsTbsZliafQUUVTixokVMX4buhh8lMa5yA
caYMqsChKzXpH+r4p/lD7TNf+QK7Lh3FOeZWgMB9m0QVdks/EKyNbipwNU9cqJ4de/EiwmIRVuqB
sO3g9Yd4kDTtNwsvTBd+aDJi+VinQm78DzlcBM2AplT6a7SMd5PDqIdQQj2EcjebT+z3swdJf0xo
IKz7i4ZRF92OlEuJy/NL7p9KVDezZg1zBEfvsek53eTUpQgGlNYAb6WiI9W5Rf8NN0nOQiVTg/AN
dCWHsJuyOLHx7AnixIoybAV3PP9QAgJHkO1bnY922gpVjZUhjiZlbFeLLig2Gx+IhVbGZE3DFyVJ
hGMGs3QiklDtEMoo3JcKpOUNTjPtjk/su96AUhPftCFOpTf5HtRxNNIcmgQS8BQK42bGSTPLo6Nt
J8dn4hzQ+REXNNE+yreAwAIpqaTXCUErX1gWCL3bXWD0rquZUQO2tWrYD1OH4hR8OHkwf2RidTuE
wIV6AhPdftm+MkPQaLXn+s5zK6kdP54fAl6JPphjhlS2JmHh4qQuxp9HA6c4Ayt7Cs52UFtK69As
AIb/liSeojpxvJkujROE747U3bwMFjBV8btXWTkMnKw3D2ANg7M9qlwERpjv684wrDyjgajKYC/F
eONckp3zbH2mth6uYvVTTzw4O9CEGszkOcXKeRbPWXGC0qhOIpvcLJSrqfrL/nwIsYuAdUDzrVaf
fpobvqLp0EG61XQvo3DbJI7sIyYoLVUxdPtWJjV7KDrMiZYW6sqbV0FnwnoJaf0ZxJuFlSM5SVPR
BhZqIaIbVTZ8ZTvabeIENQjqcNp7DzTxS32FpkkQJqVQ9Pw6ZfsKJogXy4xOUm7S2nQhl6YtWOCS
5nR4oGIbrwb7RAkIMpR7DIv1KH525HdGsCJmFDGXYS5Pzqhtwp0Zk5BVVdzO4JffQzUiUyIk2HP3
pL/m+HFbY27wAKcaQYX69wIvKfDyGLVIbAx8sZYc5cwU9BXUcHCnILMJGhqA9JF9n9GKmP0lIVmS
I+JgHgaxxpmo7HkoDSOSC+2wU58qYS4OCtki75MhFwT5/du8rv66JDAMwyWOqLlnfdUpvcC+hfrt
6vujccxhwqCxbuIsgyJz750aLLza08Vo5bakMuWmH9gp2cZlEGF6wRalLE4fOd9Iprujc0JVF93P
9yJoHP3tC9Ur9Fu4zSPp9ZVSQNroNzEe1L1b3izO2JEaHOGpv4OMTNAkh3YZrm+dmb533oJDe39P
kEixFaxXI02sT0WqwA/REhstCaXbdZzZblfSwdFtDI0rrOQcP9kCXvndyQ5p+eZxQ4W+jH23A2Lg
59uPb0EkHBpDXPK7RaQ8E/7iKLDyktXTE/BvX9dv+aggj6BubMUPojC70qeDx+iGk+Wpsrf44x3e
lLwx/wdNR3JCWf95pX+tNghqTsWt/xfuVf3qZw0U+LTwKsBrl95O5GKpNAdgtpgOVjVhU2k2iEOV
IBidzdTC9TG+fYBFBMLfWOfzobh2OBeE2bzukpbEBQKXmJtnD+3/Nrvq7zScppkSR00TPfqMqHk5
15PR+Ekff8DI6yl3dQhDLRl2Zcv1QZB9cK97mCO5xV0+EfDDlZgvpkXW08ZcjW+yegFFys5kIDeJ
agj+NDq1nE3Sw3yp3ib3yYHuPUnqjo98tJgv1bs/O/xcwQ1N+HiBYDd0Si2XRqPbAHKldlqeT76z
ADh50dHfSf68dfVuv0keXTpPW1qWGZaM10xPESv0CbKK9aBH9u8os1SrKMGFmUzS66HfFdDzZv7c
h0q8f5FuOUSIZ4k39me31Hn6pFbClb4517BO8EmyFKB5zzwZRSZVtTAuqeDQDS3MBsz9ALfvZdLr
obTAvWknaLpRsewBy2jPhB8VhDsWBGtZZq7wWt0AXfF+fVK6lNc1C/agmhfzdHBYMSVJstgsCkbZ
bwmYhY6YC7QmYpOiUMDB+MPY6itBaY2Qhm2hUiIo88gD7HvWIaW9Sb2JExNzB4WtUW2Tz4BKLc1f
xYZjzqIyGW8tHi/gwOnYMpLcBG2KGjh/nqYAhF2ZB8E2VKSoihJTzvFYRUtssvsT4TC+uetj3VwS
VIB8mARCyWCNgrvVN9oNeh5T/SnPVRD7JnCKP16UvQ5HVwndqhqFpVjiVUiaH80j0Vk+GTnqIvP7
T7yHsPIx+d63xb6L3JEjeEPIJdac4ASGNJLk3XUCLvBsHIirdC9+wJKB53OIhgecrBfIL/q2YeNC
4n0/ut9N8O2SmZN7PwS/VRRQs46JN6GhEqQrpjjbck8UDBLO+LZcAc8Vln+p5NGglnqH3FuhNrRW
UgvJ9d7tidDFBk7RIuGJkUydQrtkdIdFG8e/0N3E3MUDj6ExIEjRGNQCZKppHgnmJF0lGoXbXlIR
U51v10nNFmVyd7lBZiQ7qw9cJr0F2kwYIX7bhQlR8B+Wj8JqqHQXZ1tPp1gBetV/UlAOUEDD+CAL
8KRokqIc15ywnx6rdv2AexEyFywvByAgD4LdaXT78Jj0bns59qRGcz0FnNt2Y9EsGURMBny701eX
OewRhhg5o33q8FnIlFM7U1UFbplh3NZznBpbGxRzCzbkYjdu3Wwz20M+Bg/5ZympZ+dWXmM0UsUF
EvMXX4BZI9OcLYNGCtO1IV1sudUKJpQD14xinUyGotMMhuSRSccRTIBaNSJp75In0Lzybmh4so4H
jKe3Ls54/3nbYnW8ckaNSo7pxYLIMMFZJF0MTzzOCl3G9VyhbgOXACzhIl+U/WZ0hqWN/UI2c0Gl
vSdOGbgy32I+PKfcAYf7OCByj5f0glIW+h1vVV0ixFDbRXBZD2OE9J0Ipj/hyba6rDC/6wniKd04
hNtcmdCu1dmKzAFtH6HWq0XLoyqwYh07yJ69PeA1q6222rezaDTJDcSicZtczCEKkwcsZF3PIxi5
wdGm/4SrKuU7aJM/leQOQ0TS3jssvjBRnVtenuZxLb0O40oHJ5Zrct90KVLMl2E5PWwScNMpT7Wx
6wSFUbluEzCDWwIBPFcLdgh2Dq4n82Dy2M7TVoDGBOAfFrTePJwGWsC8jBAdxNkX/kkiaXMJw57f
RFJ/Qu9XeH3gChBCEfRYtVd4/YuYaPaMB8wIKQeECCJ6PvTDrPzAeMPt4bos73rqT4kM0bKHXqN0
7oUYO8e24ZR9Vuu082mNlGhzGPnLR8+hOuMlrU1nbHj9saf1ONlA77UERXqTNnrQHmDU4Da0VsOX
MOsKjdxRQ3Aqdfke3kKjPbDl+mP027qR8cR/sxISb6/Akss4eW63TAtXFXDkgNTyDPCTZImpCgpj
6WC14z12cotmeVnJZMIE58jakPCNfcdU+WEoFt5dEGT4KWqrnfXxNlbdVOY6I5Js6PysT88Zxi8/
lGcyXtyAo7qkgaOqy44CzqrJb3o6XwPq4DxkfOGpoPY8dFc/TpPX3US6iUYxWocEoobXg4TwtOeE
52b/IrkNuIet0QnQYDlOJgXv69F8CcEemvlT/VNaVGMFwdc6duVLkZhELlh1dk6y1KtuC6KF4tdO
yQWpOqK+MQrY2XXz10JgOAyCE2pzmXFIlyOkXE6XNxstd1eU2LE7W8EvzIH85K4GW7p80hYnbUqc
hKoYv1W/C8GIGi7PE+m5s6SAODk3efPeCFjlaBCFl0xOfgHYR50v6jF9+8AUK+TeEuN3lJo2PQbx
QTMKTafv2JszhgS8U5m0xCTA4yVHM162iX5heLkEvzIJzzMtIPEHURe2HENI+DL9qslOyPyh0O1S
j9yhro9BD2zu+5EWIe7G6Vjf8cMWMCVZe8cErrOxzNsT4Ww4eRLh+9nMwv92GPV0qKmHLVqN3YhK
Wn7BQWIfp3LGqtai34PoO9X50ClyJaWv2CjdDi+RhRh7cAlZlqLELbXWL6mvs9rm2O6ayuv0s6iL
fHL2PpYra+VYTbJK8l4o4U58SPiAhXVDF1vj51EXbG4R/Sr/aJj4GwTGLs74N+f/4ZuOy7AWSDdB
fnHOKOaeJVLae9R1adT2i1zfuxy8p4pf2LUCIvTyXnGTkGTu3FKT4bmR3UK6WZri3fyAddmvy8B8
69Yo1+2SuKHnf4SO4CpZJkbu7zAuGd5ZZqqtjfOZObW5YrlEqwEzAmqgSZjdEVV/mNodlcp8PiVc
g7kCsflodkjSkgAPCQkWIUR8BeCzOJT8tE7dhZI+3lTx5OrmZ+gAQPlbAGaTwRaSSYi4lj8YlyYO
VEroSTvr/r6VrdUJNQwLJZIHGcISX0yn9toyIjKJjfklh1FnuY0YUdxQYC1VybAdqTLHcNpPhLZa
UA/sPDQJgJy6h2vqEBN2jmVscLFTmL/Rqt3nK7pvG4C6EvZ8vSwjK46bMtWNSfi1LJ4bZuqpPZ2m
vIa/TrPnfUqFkCyhZVRGV2r0uxt5neltyHelrIDu6GTLakLjb4eF0CmH+wd2VI3lzf7L/d8gilEj
x2ukY///Tr0pTSiY2IUCAGLklKaWO1dteIRo21KF/ub1hTbwhcXq0Ao4BvuV5s1zLUUNgFDg0d24
UI8SmmNYITA6xBxb+1Dpz+6JM+lyK3GMlB6IgsDNNIXV9YhIcKE1mZZCkLWSSCGQq56yIYv0151y
ajhEoeXRInXdmQlJpse8YAJ7KAVlK+wPxngjym8AbRIqEOo0nq3y1L6InHk71fCHFVFr76unP1Ey
BFwzf50qZBzjl49zMWdQZ4qXmMdVSgENxZK23OpwiRb0zmOVjwK+Ofmdcj/7GJJcTUfnRpiwrQx1
iI3tOg6q2x+r1PIX/mMohI9G/6uBaCQKNMFYx9Jn86uB31j/ARNPE2Mfu8R0NuRXmtt4R2x4ZCVC
YDpGe04+yI4RfpWrFxbqDyx8JkQrNyPkKEx55oaXkLpWQZXTCEFpynslAzBWDJqUwHsay4yTRFdg
uVwhgF+aQSEwNlMWFBsdpvP7o7GOvBHP3bxptzlwmd10Vcp0mHQXXRKfoMt6k2wDIPOvTm14uRS9
MnzuWq5Bv3hYteHrENNEGz7UPq9Z+AkB+W322oUHt/5IOgx6S0MQvy3uGQbttFZuitsv2RAuOF5G
VCPEs7d9zqdKEZD8vvzLh4Mdpp3nzZQVijpPqWiZjxiiARIyk9qdvGe0Mxe0OJsH5fGOMkJzuATv
9v7+dfk0LAUEY69iY7zGdBP8rxx/g679DgslfKaRts9XQLZJ2ECsWIhYflq8Y74MklA9sso38rHO
bfHXrnSW7AQyzO9L35PV1v3X8n+zmRrKp8Qa2rUzaFPlOADOuKoojU0dgjLFY6kKGAW2K9ZAuzat
DQcWUaq1VqDyjlgLJYEzM4gVl1Zr6VkIkbOl9n95b6erlCMGqbuT+UxanX0YbUuTRdpmkJerLonr
fQb1TF0P18Eop2x/OIO4QlCECCV1Ly411BcBJE9/jQ+aEDvxjP5rHBYEJ+2Gye4zwXZRw752tlcz
cDcPsY4xSfCiat1R02qQaxoihApVL2jlmaxfem5kIQ7QhA7yYZIBdStUYOhZI9/hyNe1Si/LDquo
O7O39r0JZUylQSLmHUhreKbHJyAziwXhXP9DSfXBWesQUEJ8Uy682puIWuKZ9heCfgsvij4oeqwI
JD5FSKjg5Xi71cprXKlUVxBo6ZYVzzowuywYtVEewINA5zJ1p4P8ethEk8/EkOfh13mTzATejgz+
PWoFo0GCnNgC4TXcMWoDj3smvaAUhdhYj414cIpNCz2ios9Dyp8Q2WPqDt46U9/uoJT9kAjNsqLa
vbRZjRNnhkCg2BYHrE/bWAQNGbhRbQAwmfiM/0mJyxYOcs/4g00RDGjh8zeib4R1iWpjj6r7N4JC
S1YB9bQdhylO06O844gPXdqH6PVKe13I/o2ivHhEkEYjDPWoys+JH+/I7omrRXh+MTCBr8bNVZYH
j1PF4Lm33Pwzey2PUncnzlibl74kwIPqONeCtf757cSx89bzgfbo+hPHPKNQKJh5vgCe9a1mYrFy
kogWOLWR6BfUsmi2Vt/qzyYZS2GjaCgta3K0XyDeyrEZkXHILGXUW1Wak7yp+lwR9pP79s1hJsjd
rwQuDJn0PAbonFUWqBz6HBljCJ9+2WA8m9pabuwPxsVWSHVIi1n7ZvMOLwuqK0UY5Gn/qaDy/mI+
4A4IGp3jJXpASyvLc9LAguySBXtR0IHDembI2nW62FQrvJuKiwebGuk5n3L3ZeTCXOaLLUKcN8Rv
Zwd06+dKAGWDcvjMbl6RqGZUWjx2JTXmNq+Z6hlG5tCYwM5LJnzkm5EJ6cXBZhKHS/rEdZfbYfab
UanbJfNpfOz0rPTV4WDJ36NVcXhdYG0UgIbwcDkIUpNozis/41D+Cns4UyIXe2NIvi+ZuMlkze7P
S+BPnHPjldsODGsN1zY9bayPnuKbPNw5eHTtdqvOLWYz6D6qM1uwfnzU+t2b8wch4tbVfV9Ia5RL
vD6vTOcZKFqkd0zPA208vMaZlpV2OYATCNxL3An7BDDYC9MzOYJEzEKy1kMzxs4R6jh94Co65EvS
qYMGXtGPko4IwY4WI3yJCuMvPcmoKOJQ/+hClvMsNjh4xJb1qmVyiknGIzgAmCyTMpUXe42gz1my
DOOXZPkVqrOA9mrOiJH0ZO59aWuZyPiGFCWDNlxl9Oi35H8zsSMJhWlkftmLPXtmFMXw8fs4w+jw
r2kkbaTVDG/zNs8Vvg0r2O3WD0QzUC2dqwLErSzgqK+t0jraJaz29RAyc0gqM9oVjQotdsOf4M9+
/TyF3456zjNCHLU4gKb05FJKSEneobn72GSfw5QrZtm2R47r7dhNmLEMbkle/J6yzymyvmnlyI9D
gyjNaiOfnl8YTiMrG0gbozxAM6t5khO0hd1ZZLtWquoxXcAX5pzo/2HXgpibAsicVHagG8+zgIhU
2O9tLzH5l68R/w2m/3EsjqVpHzqZRTAJrxhHV5Obbn3OUTZzhb2CGsM/opj558VJkFnGOr1NbqWC
WgwGmH7uCEyTBbQrKLj1SddPaOiUTWw2SXB5w7zj1AKsZKUTIxw5t90t1l8LcoK/cVZj5BHZPoyz
pdxP6hVkEscYjdmWxuzFdP0L3UxIrwktp8peCWosWsv8JZT1SrG3AUoDmHKCSBIsKFlC55RKGmtN
1NeHB6QW0UkvRwEmagw4Oi4ZZiueTmnN2ApY7PQG5zhbYEnFJ6rybg6hlZv83pryV53rplgaNKfn
FAXQGrCTbUzD9221MKLukXWZy2cJmD8OxaBdaGoHk86IETkovzMc/r/kquDHJahOc2nYQqL3lYBA
iB4C/UZjdttWuXy5rDCj4wIhl/KNQnB0k8S3bWwWjcEbXiW4uUdntj//vMBRgp/sbfOpnChvtlxQ
ZXrOzdN3gMyEPTz/de/o0ap+svaXf2LVv440rV7nneoGgniU+egD36kNdqQNcnJAMx1dxUidkjx3
8s4UwXCTv/fvyO3GT84LyBaSONHip6cAYND6Yjaj1dxVAEi8X2HdbPzjWgWwKwCkuzRphyjsW69d
9LAT7Tk+BSw9e8po6lmBqnttC44OVlPpCZtK1J1OtunlCUWem7lBoXBvAGLzyrVIeRJklsSlUftv
J372PxKcJyBpvJaaqkZ1O4xfIdXaZD642FbKlJnGt8X0+MsSYsqA4/wdArdrSx3xEPFLO+GCCfsp
mCTXHCTbQXrQACnbywiiDPjsCip76qCneoOmFVjBXv9dT7Zb/zKymUvGqmVAc86Dyese2D8w7J53
VljbOri9gAXiMBG2CJQF3PQeMk4AA3bYH7vfCtvmSvl+b5nqqAbcWmw5HK7krY6ornXkPDlkmtJd
P9yxJLtxxtF8Lnv/Wx+rajCCNNDcxMOieFbZGkXPVu4Hco7brKpHqCi9bR9l2R9WYZ5KOWUMr7an
OsOnZ+fi/QuMiZTEL6rw8uVLjMLaJD9SYD7YtzD1ewPa8tGJAaV0MNIOc0zfOUJcYJg9MSm8hhYg
v74iyF1/ye7pdz0wokGvzv1pvJK3K2KAYGq849XBbp7HxsMiuw9nsASR9GEz1y3v1zg9PdPtU/OK
j24x5VFiv2iYYPXmJ/x81le6ZbNgots55C4xZtBm3nSWvNkk20u7WSbjejnSzfClOdR9W+EDC/31
T9wpFoOq2v1/czDEJKJngQaoEWk6/h6Tr7+0RusbCgH8XjqtAec7fucZbu89/zVWj1gIRy5XUrDC
5TBgySj1AYMats/VoCCLVyIFm1nW2kTzvNSv8x4cVT45ovqacOkFZEVT4BS9RqiDGizMlO1Vni/r
Maacr291P+XXksTPr+qz4Bv2BF8oXyeBnINJGzPHLSjOk+h9wBaafZ/wHVJWj/bPNx3HH5DbnihP
neP4vRuwUvHjjNvoGEsOVuOTa+CZWbxqc67gzRUnNE3MzIKjWmRrBsbTO4ZO5QlLMb01bmMOyyHB
9QSBp3BNhorzQy3ubuksvCP3GWeAEXAUWFs9njouPDTcISy+6MhBkqisinMCLbvhiVlrnpKHIvRo
NC8X3uv5b2xJ1oinfs7KjvIsoLDplFnrKkMu3FeR2y0e8KJobvOr5a5CvnKlhMsf85sIgqS68NF/
CKyuSMOVYU80PXFR5l80eqrWI8jtw2wIRROa3b2wF9fHyCC/1Y3Uwrlhi9mzzn3A4CQDETYC+HZs
7MQGxcw9Vkb2FYUX7JisgKVEe4+WuuwDpwjehiSb+YZ/z+ciPJEUQFYDkMLNf6fMhVr+MazvYdZX
tNbXyqf2HdjqIyEJ4Nqso4+vB6QQJRNWDooAZ3PFFluBNrDNrJ+P29xT9Zqps7BSDnOMvF1Q59WT
D/stBQF7HA/xMLkLyqE24Nyib1qQOB/L1wyCGX3naA2JeYwuRTafEY97nrFDHEbGBBRnjygoZRGq
bpOcDAAAKY9TTP5K4UUmVJ+FT1Sincuo5am+BZZonjtz1+R3wo/+7Y7EtRu0/i9+QTvYfPzcb14I
aCoLBX4ZRGCrCKC178y483+bm9JG4pQfATCznj4HH+xWBBq7884sBflWNkBV3kh3ZVnxhga+T2Le
R1ssSjSclj2Nw2QS4PGWr375sLVuJQQUZXKVGti5+sk46r/AI6R3n7sfR7bbsNSVDwB/m/TNgM4S
7Biys1a5dblZBhtNJLqU1XxPN2COhiQLqupwSeWMzYXIoDp5MvVZgil9FpkvS8VwgABQjbKZPmAB
bC/UopkeU+f1ORSouPFdRsRN/GQkBOYtID3y+x3uBcwAepd2/vB2zOcy0XbaDW3cBbByKnVs2JsT
SPzE2h77VnjVSUbSR1e8eNIvKuoKwLPZFmMre77YusMhqxaRuV+lU1BUt3Temni0UpykYZN/BLI3
2usjGrxhCByK/sP5YVMCtUwOZszrBt22sM9zhmYmAlfRieyQ8WLqY/dfLSD496SIW+Cv2/bUluFK
60h8gBAmSV2rPXUTrBwsagpch4w/eZbKy/1e1w5XOAzeA55I7aauw0mO0MPHvfpptLsx2R/0Vr4q
qPCiiE5mtK0KyvOVykeE0YBGMFzwTFn2QocBLb/OITAZvLGgPawrgBCRVat1ceRTopxD8f899Ef1
3kmXGbRGbC671EI3TkHrPD6CGEXnlirSz0oW0Qgt6dbp7wnkJ1cE9rdAVQOK0fMgjlnA5q1IvIrG
WlBg1em2V4tB0VYrXCbgLDk4TDZ0pJAM6VKXnO2/ct1ibwjy7oquwPwjLbXLqCIzYnXz01zYrTor
PJktmpzkWgazs2QZoISVNAz0H6kOIja4ke1LJY6mGwrUL6GuxpUsPanqCsErl2iHRlsa3QPgg63t
6plILAcofmiAXogcme6YamIBP8Sd0nL7ywV/afMaaUIWx50BMoeRDpRe75dQ1kVBJY9H0nRweNcG
5lnacmc48c1x0EHHgHIA7aeWMlZ8/Nz6R2/9A8w49PwpnKGa/8Th/xECJjhTgan8Bo8NBOdhPZhv
E2xrRT8WWIwEIa9kcpw40lcU40es414bQ9nYARwCQsREAm8+yS4Lj2uEZ/MTNCmKCMekSTMcFQ+H
0m8ynVgTs3LnOnQaLX8yoxkAj3z/tsgUvuclAHT4laBe/c3e0pa/Babz5u7ZBp+WZi7Cp25ENHLp
8L7MY7g7nvyPQMZbeNEyZLCV0A5xFg5EtjnCac3LKE1NkH4XzUaNPK0LRnoQMuMuU1n/pxfx4qjc
TdaZezeOe7rqod12+qE2YmZiYDnajaP/mrsXlwOC/vRLvJSkjlyI/BshNbqWtxX9/kRLcL7Z3+e1
8NtGAv/N59Zp6kxPWblW66vqpLjle4a9FbY/GfNWIaadrpB9kT1FJjOxkeD9Q79QLutWHzeETtYx
n6Zl0BlIL9Fkd1NWsdF3ir5KTpPYpy/wczTRHaOBOrb3482UevnPw4kBsQP/wD6NhNfzsr1d/q/N
bMnT6nBlPv/f7p4k8xvDa70dOMZhVWnROyPQgFz0nSXprF1tb6zIxC+sf1k+6zkZmY00ekKj80Qa
bLhYUCPnzOc/nfHjt92Xrr+6gPbfaAi5Hd6SLWDZGlEFAU8hXWE9jXzy/l8VmyOlLaZK6ftMeqUl
vQZkeESZJAHUT1wi4sVI6Mz34l12jQ7vRWb6iF+4SH9W5A1ILneqTlPyYwetDMzz/CYPWAwFI3S5
8y1+dNzDFmO6BxNZMmHL0L5i8z6xEWuXB8aO3erhon+JKQwO8aPtoiN6igE2ZT5tTldeRgGluZOm
g+7dDEOymY/7X11k/VriF5xlHjDJTiK1/udUMa+c4RXfGsRteWJ6HFl0iEmiuENXDS8uBNdc/zbH
E+bsvU495j3xdXIZ5DyU5PvrFDlAH992oQZma0cjdX65w2S69+//O41LDIeOqWEfR7RFHS0naSnZ
q9Z92WCZnj1wpKIk/wtd961hKkQPEz44Ne3Lzg85AC3F0lAmunKHgzh9zgSm+FvOOxrQ//OBTg1V
LM5wBvUZxgN/mkVmrWunFB011DKZ1rRNoy7ss8JIxaRvHzmXeiLdhUFvGB/2MKt2ExMoYGdGAbvZ
w+epF4yg7DGyyiKDRE5rg7N/ZyACMH4eqebKs7foQINz1Ie5TZsTVgBeLbqAHDE+VNVYcriyAY8I
+DHDDGcfYmjz8l5KGUr419nqy/WMKZVPy00j7UOrIqoNg4MiIO4a9idIHpRtLlKZ3aITZlGawd1Y
uz9DkHA3xfUd407Z63eV6UCNFlASwTFtBbUnvlte+U3EsRapmrJsuqtEjy+k9Dhb1CItwpl9i2hv
1/0Id619Dz9LP+fenkq9DkDspdHQiu2LLci++QqAM+yD9YOQElRNiXl/aq9/KHO7pGQJ/3G+9CHw
oE9U07s76XDgaD5S83papkXeRzUZoW8wca53DzTvaRN/31DYAwjeA1R4aZnOg58iCA8bZAMNleXZ
7i8fup3BKva5bXWn2F/wEPjf58vZmuj5SHwPsBce8d+3NWnivdNdljBKRUfWHznMGe/1b2m1ORMI
sn66piBN4dO/mZxwjvG3Mf7oeKuEiMWHNj1huYxW5HaKdx0UeesAUd+k/njg9llyXe5X2uNpEDOy
lXylTKuFSYSYk6YGw0Iz3YzpoNBSkHNRgOYYr4A2p6AUQpyvUYBuKtboNVglajFWhWPnUEfN2d1w
C6K/C6a4P27wuFZIOeypfKnKwqoGEcQR5EH3/drUe21h1lyhPopzVPOR0ANuOaujLFqO4uncIUc6
CqxUs6P90KiTKcUPcoVWKdflhDFHmlS3koJsxfXCKfmrxd+6euwk/2yYZ0ejZtZBiLKXZkCujER1
UQkY700YgJ7rL8wdWyY0o59cmo5EKPLIzL7Pqm3xikitHcpc7wIf3YtmA18uO98Sr/88ZL7mj3ex
RbOtujZZVdvghEHWQ7fjBwtyZKBOjnKi17fpQi4IvOfoI0GCXPuC63ADUO0kKkrkSplSBZ76sOjR
fJp/bdIZUCDqhALCfbeRlUy+W8mvAY/et0Ji3rnbjknX9TxYoQqRl3w87FFymWOqM2+tMC4ZGete
f+ckDZzX72EARBZ6i6Yyl9WZ6xQu/s01yUxoASH3RGIAtw3w/trOjffmyk7/koRw1j/dmrIi5Kew
kwCRtzWcudsU00thdUEA9AtDLRk5uaGTAws720r/EAF8v86ML0GA0F95Af2m+KMdiVSV+vbqL0vr
yrWoLSq45wHN2dkUwYRWDVp238bfibViKtuSWg64ie8gDqWNu+HBLNUDoJwFMmcCH5Spl8yHhPBh
FlKnqiz3iBfAEecEAJV3zqbr5YPU/hT34qnWjEhvhcO7P3f+a8DHjhFn5c+0H4f9Nj1tlumgcYUo
YvHuSd+OQzUU7EfjjhgzNb1WmHfAsL1CHn8sDG9xDoBx67xwinE/O2ykiEFTMMSt4Yow5V9EwFac
Ke5xZs12QDG5NUbpBj9A3f6aWBwLLoGmPUGp7B7Xb6Rgctsa4AgZe8aahwrV7v+wscDKWb7Psroy
U0DzZqhpWluFkurFumUlc+VInfrAMPjCtMKrJ/1z31QbB1ZVKsqh5kKAU3c86syOGBOiED3FxSx7
J43RXeoTQgz7fE/lOiBkSqAjbc4z20hzu9onR4bWWMjheSRRgbPQZjuYwBiM2d5nwSAFlbv4Vobm
xWqYLCkBIlONv/RA+rpmlEqnSc4Cc/Z+FehNHsdMSmXdaLTZTPzLrA1hKEL8j8cyPPubxFyeUMph
1Q6yNEAHbkaRea3QQFoHV3+JTU3qdtFrqHjEdOQzXBQesoQf1RV1Y5lbprnKXmYHVc7gnQMLwCBP
tB+dD7GI/cD5xdU0jgkkcdK3A+eqdOn1jfjfb6DinaD0Hr2mH5sfFwwPWzelf9nQVShN2Yg0Ah23
2ukF9Usg6ZXxcWFypUy4KI1mW/O541ZOfOIvET7y1VYeYFuap2GCTLDDzcMDbidaw4Hk03AYj7Or
0CWoPJYAdz4Lir3HZ3/Wq/pn9e/DCP9qA8uEXH2Km3mfmvXsV5cDi6saF+NH5vrm5J6U6OJhIdOg
oN9XGsigY9ykzgnbZKx0fUCyQb1BO+hSZrzcBmUZtDDRB/Q53ZgPc/SkBUt/ek0Gq9sDTyMMjS11
eZ9nCEBegI0IoxkQvgcjVGfkoBnufI2TkUGZo29nr3xmKbWOWiwGls2ype972g7aAFaqp4SY/qKK
y6dXRH6YPEvHP6BRIT3/wEp8J6fNoCuPUMkVJPuhH1LA8rEcdHyeqrHyLxsh1WmVAsfSfPVk0MLf
4H/1YIxwK3eqMoGc2QdWPo7duFU+C3NmassTOpcW2kYcxYYBm1S20UKCLxs1oMr6D+ik+maO+dAM
1UGcPdbeQv+BDmv2i24NkR1lB3TUwjLw586KOmahZFrx9635mDydizKGt2jJQfM4NpqqBqrGui3z
pcinKJRedlYNGOtyCKPTEFBW9PudnYFgRW988qy4xZ3p6MCSicRGaHVsI5k0QGnUpbItz0hBY0ZV
D47m8g5vuR5+q3I0kABKrds2iTHjnGiEoMnTQdW9GQ+Bg23y2oaa/BjQXPoyNMM4kRwEfaoW/xet
eKZ4B6IwnFObdJd4nP+BGSV9A8d7Y9KK+rN/izBAbJuvAd9atkZcULi2WnIfjWrRtKA6LzaObhnX
wR7nRUSAcox0No7s6zB12Ajc5Z1LaD+C9sCsKG/NX9LO9pA1UXokaQtyyCFlqrqgK4JaQZC9qCFL
WlVmPNXy6PxEKp2JX7X+v0UbbOajBnMrQZN9xquBrZIrl+b2UCaQLdOdc/HELXO1ZYG9R68QSpjh
FdgbowI1YeyeokZVmBwhHvg+7/EtNAfUtd58w3+87+fBmBVgPGes6RPP4CBFLPHRH7Pm8962k+QH
jXaULP/sHzbuEJV1bcl9sUavI0bBmp6kIzoh124b7vEJaALJFc6aXA0g3ncI8Apy5uRvuWnsAita
DX6xQm9Iw96iJGGgIvJQzxmn8IcxZmWHPGSI7/QkeAYuASTAkkQjVB3K218VNOjZQ17UoR36Fmfx
TYauon49wl40EBalvHr2v5QjOTprq9wCVQqE8PfKSxgpr5GpI4n9o5M4TW9w7eIbKRzt4wEqWebm
0D9vm4KhAMz6nW7bq5BCFu9zIGLYxqAN3xvq+MGRLM61tvepKjwMmp0TqCLm9QSjG7pOy4x8pSMm
edHG5XNSJP5LWBFtpB5ni8viIIJhFOyUu8M38y/VWEsX6pIfE/qxs0ACFhFpMaLW46+XUg4Gy+Di
KCCMY+U2JOKf2V3CaQt6ln0glSxq3pTtvbZKggCx6lTedMbnbvBczLfac96QABqfUwa4HnYIbrZH
OBWBQp5ADJ6+vbVmRfs8Dqxtmke0ardwpm0wl6OBvmWXwvdL/mkNcAekm+juXA1+fKQbn9kwfKU+
tGceRHORLGisjYuo00Ssp00E5wRp/xWBcAx0o8eSXS5PppIly0yVaXKl9ehIKGtFBazQkp1G40Fy
cYF6Dx4Uqs0ZBK7RRVqOinUk2MPOVenXH+oF1e7RpmKUs3iGAsRbHqhRMh7NsRLnKcdSQK3Fh/Bu
keP3xjKSjNuozlsimr0lTbBzjMbLGNKr1KPb7MWofkFz25pWIhUSe+nO2agYtHlT7RzRSH4G1lmK
aXdnnZ2B0He4swu0k0rvwHjArTB5q3P8M0io2Vjq2rnvZ6K85cj/3RSCJkkO6bQ9C3Xe0KaswSq6
EFrrojAMuXEq4qpjWldDZVNBBNxkQNCjnWJn6dJ731f6LnYS8lgcwuF6gLx88enzkvIWSTu5J/g6
Ihs7RkO3CTkAVyW9NCSw9niIbS2Q4jighCRnWTTXUWiW4B79rFHuQIGdRHTkbrEVgV0zsRHQ+ALa
sb1XoBtWMvwaFmojZYvh1T/XC6Sqp3PKWp9es5hnYfU+T5lJJJRnpyhb7ASLU2VMk4Y6bAsk9fDb
clXPSnhKB2D+fiEz4jrAIFO9O9+GU2Vulc28fVy0wnX9yB8GBwuKwe9qcuG7kFqa0Qi0bdNnjwJh
vNUTo+XSN0VHBUEg+w+WJL5QLuOEdyO47xnCoT5Zad9+7QS3PbSkZmxKeuifBsJeGinhIwrEm92h
l/KCKWAyPX36FhbF8sYd5AlaZBg8jVv4xkfCsF8DlLKRupTw6DQDl9dsOmN/S0nrmywJQLQ0hPQN
INgYkbTsOxWLLcjqKJF7358IbqzTTFjACaetFF0hQLXg5VfG2vzIHM/x6IpYAjt2dUT4mmbukwne
/GIzhocoLTb6ENQsmZ0I+SG3AHdYfLb6zFdYkGzT1d16NTt7aNphcOuxD6retTGCs2iGbrULHDM7
tZbLbsE+2c10gQ2AtprwIkXxFGt+SitHop6z25YM6gz1OPeIY/xSr3NfiKvw8mHrM3tckbfzXaSm
nQXQgRy+TTPweGt8MkTBLAiaF++Z7YQIPpqgaUGx1/mUFsypr7UKmcGVfSMN/9pZIr8t5dMjzkXJ
s15ad7+EGmK4f8boC1lN3FeFBmEwuS88jxhsp4MvPu9yq8vGqynfMQyDyj5nbC4EHjPY+O60haV5
52ne8A0ssSz3sv4RXidQGNij0QH8AVCp+hAHMpQwVo6bqrL7F5rxMdURv/9Poele2ALE8EE9UuD+
QtkMpBI4zs0qw08Q6go4Fj7OcmBxT8uSaSHljtcOuaYm3OIo4Ey9U4BDDepD9mDIXv37d/RLrCpJ
/J2ounQEKT2PJVWPTxNoMT2w4BgMRiwSxqxzaLUENRMi/MdjdjfFF/NDGOqWvgMj0GyvUPHaf4U2
P/vG2/SMBd05EUe8dzXgaLdL6uvneZ/IkU/PthhmqxVb+79xW4FCZwUH8is2It+gfbtsbBjWi12w
9MseFkvzlXUQlNXLIHJt7PfrnCvE//Cs4mQC+J8gTN5fH5S6DF0J6oQ9GIwIh0WVbXiXzunXQoJZ
kc1HayOjK+x0aC2nKztwLh6ihF7SaNlwE+GG6fHZ8fRs8GYwSKbv6u7pjg3BZJOPLZqu+aM5iG1U
fb2v7Hcz0ywiidslsdluqyDZvgKwxpkMNwBZFlqgbLmCaaJ05V4z/Xatiqtyuj+kdffCOK73BrNO
3ksL3U+F1KgG3c6xbFYWr9u78dUPcDaSVJUmPWVJKC0aKEOpBgAts/nMnae9Wq7KeFfzZgHhp3qF
6Jl3qff3N5ZDOZVbOATIipEI90BL6OVwBJkcMY7LT6wbdNMgdosHCrWFC48qztgPHdjQPq1+IEtO
v4XSsM1qOle9vbGw+y8Elxmm+FgFskmSh7szcs5lu0FWegruqOoBXipvcmAhRv3y7KyYU7Gta1gf
ipE08tkCEqafB1YS+DKroqoy0tYIATHccejXzXQwg9QGktJFTuiYhNzYy1cmc7p+ArGMkjQMVsZ+
9zqY0GSuB2dBWK6emor4ik0lExek4h2Zoix14G9OItwlRdTaER15XpPdBtACElxjwtqnSbq1HIRd
Sq8KAJz29PzrVr4CLT0T2k9dv1sOgC2/bOjJEwAW29ctrp0Fru8opZLGQ+EPrcvZQAKPwmoJK6oA
b+zFWcEgniQfcrtrwTamFLmmWPNT9yMENNbNg5x+q9dLZJ13oRNsL29MNU5jUapTkkKWqGLZLf54
QBg5zH+dkS9JGBabKAysFIpuIm7U66sO2CcmsSe32HgPxUvJD02DzVyPmSjmdBKA73++3RFkrWGN
NXtuhqC53ZRr2PU+P13kpVUKTaDDOgG2xAd0XokD8vjz5KUXA9b1YUsR/sfA/kUFAFCf2uYTBOTl
bs9NYkw52a0fcyk6+fW+5zFcY+62ENMIVPS+/JCqZhwzHjWK1xRUUvUyrlbvW2RG5REu8h/5/24P
YCsDBdMTTjszj8usIpI0TpwnMW14qV8WdnLGKin5ULLKftqL23NQ2gn+BTxOnjznggct9dK/ykEc
vjgLseenU9cAFgrCWIAyGX9IgoRJr4TD1JGxqWAtcb4e+x/r0FKPrMgGUfxxbNfLwCGxwAU79M8l
/NQPDlg3VFYMATof12nNhrpOTtMQjEPhgUp0yopBL7G2AQS1KBBIAq8B+z4Ia0LxSz1jLhEwh3Qu
QmxgkKsZEBOPaZPii7G35pkPL/pyqVYF6EbdZWn9ziRsrkt0Ddv3PJnSNWTczlkua+H9xAXhzBK3
ryLIubsjThC1ygMiCdJYgJCIW9lxQwFfcS1gVrG+3ogXbaofKwB+kNJWnDzR+ploaT8xqEfC8VCL
uGZms+hb07rn0NP1Oxq9JQXvd93iuo5A+BhhF15bsDMiGxaQhAC0v0sIWB3Xs4CWzowDgv6z37xm
ptYiWk+NL2BzzyRTuqnBI7jRBwHupQvpCr3dM4aGlqkvOcN+6GZQH2j5/oqDS/19ZCPlOUjmE46i
oV1/BdBZHY2oPSINyWxPe+qjw3rrxVoNgNKsvU+Bggq4kUz/Yuxo13Uhcy4wkBzdiyGN+D14S3i9
A2bBvvl6sC8y7uFa2qOZZi3vB5ccRR4d0PTSLEyMS/Jf3l3qdzOAee4Niccv+7qnGc4UcTXyJj91
op/mi/HoO3tZCpdiH6/AjVe8fqsALBFg4/NVmB+iWaiUoNLzY+W6eq/c0SKTLlchCQxB3thmzHIa
LqUz4yEudgwyK+XoVSY2lrHRw9/K5WsWm/E2gwSWWE37wi54QNDyPY8ES6d7b11QVXFLw3xjLerB
I3S/hQ5gMfIncU58RlHIoY5WcvevlwZu5j0oW8OKv7cT3ZfqalZP5hl7bRdyfty0O3Pj0IumdY2i
X4xkIv5ekhicWitKsiPxdUNcjyRVQs1oGS4vJSdNYxyfjCnAVtmPz3dx19ji9hmgQF8iSyJox58d
5ph6+ZtARRJSrJbau2NzE9AmeJk4E4Zrf4RCkXjMAMLi/aZH1oKvXI9rPogcA9K5rXtac0xur0N6
powXB/JRLDz7m8VjmGbcuxGmiJpFYHa8Px1A2RipXXH5HFM46tM6Lb+Q9Tx0MM7gPki6ERTnb/YY
QzZ0rpEX8CDbwbbW7d51iTKZ2ka+cUX6WMlXKEq+Regz5ESK5dQNbD2wp6bniTU9DcwgI66fUL6V
h6tCcDEK5/tvRD1IvO7mklIeU+/9qn/HtHU2Bt+kZuMd4oBwK3FL4762NPuiguLWAi5Uc/hFcy/K
4UuWVEku2mcGFhKA8XJUFpZFWFKND/KgmLqsmzGSTellFhSyT/R3Jwfg52qXCK8BvU240y++w8z/
uJksfcu/I1RO/JpZ5j/7R7x4ZP5tXGdgNAxeDBlbXmi/0SvOqXj5BVUUWgYexZ8kMfD+Cjrko8oD
80C7X5J+wXO8IL2RI8+wACGX4l6nqvFmwcpf2LyZV+q02O16CI27hVpJY7ae6Xj13wLUSwKCgqUL
q19W8EpkqWRsc2ADB6YvE1GCgibm2Zq1hwv3lGOVD9KYjUizKZ5VoMiMqjAv1FgQuoojgVGrjJxa
z75EFCFLP0fXDtOx3cbYDAfGDP7RtPgbqicJrF7YBSP0NDI08ZMT5k6ypGFDrI1PfcajehH3POfW
7mGHzuE3VMBUFBLdOkjWHnRMKqyefE201y/54Sj+3Clh5HOAcV8uVDPxXi6suiiuYwulnBY7AZFP
minMBEjZHR/JP0Paon75BGKH6ABWF4vX8CsVoD9t5PoFXAGsj2bvZHnvx/HEHCaq6rO5HE2u6p0M
ttduYpNpXFkp0AGgKLdBWJQ3pqZ8BApbk39a/MaitzCqei+r/Eil5Oklga54aSA5GFx1j+Gn2NO7
MOHn7uMggQtmGPO64PgXOJ4dN0aolJWT0wGhBYkXt3ZhRNoig0ENZMjWWmx5HdWvX62CjsETwFJ8
3vYSHn1LkYMpj74s/t0UZnuaWM3i21ZfRCYhT9GsgSC4Y6r3eFaRe7fEMjSB+z7Z/lHk5TetAuDE
m1zQWSL/TfN/KHgrD9QQX2u0HTplsVj5vN6ze/MnxIB9l7DMS7bobc54fgFTTIChCrmKgbD2LWd8
9xzzSwE2NHEccTf/56IxSZoD01nAPskXOaE26X1jBALYScvN0sJBM19GrZSZzMctWVsB/p8nZuw9
CQfiRG9LPFEma//2WgSS6mGr514cNsu6xzpGupfkaJc4s0/BV5OTYHT4h/5VJUyj/7odwiX3Y2J9
CNaMQSvSgjLZ86s1j0aErbG8weeolsjY4jepiFt82umrxwvjTFC2DtDmDPef6tvC91QEVyJTgynH
lruZ1G9mVaG+sHxQGDqZn4inEF86SVQZQfm8ZXpGQF/TlaOQbWujVuGy0+kwF2tApxkJJ7oX67cl
3R6X2DIsmlFZsCPfRMsUs7T0mL7/wKNaYGZYfYkyG/jhOn37IF5XDAPfX4wjxpnYZ6G7pkvH8GtP
0Vb+dbpQJNPfYDeTskhc9QVYyvL2etSOLSR8qmUaqUK7HI/+fdOAsw13ZugzfaXKHDRbbHAQ7fDB
K95zeYsEAFjHga35OH0yvM4xr6n28dFsi6kOpGr5xWoTshzFBNakC3fcg7zaO7f9jZi3qJ6t0JZO
cEXffrW5FBW0NmgIbdc+HWXnEh6BU/osg84cCpZA4UDb4Hb85lYZYfwF3QMR3ONT3x1Y9QbcTlP1
GE4fIZF9wi9xw/5yvGoUyp4MhSnlHhbpmP7dHGqiqe9ENBOayRjPD3dqqvf2ubducDhKuLqVuYqe
pozUiRRNvRgIABhN278BMtFUnjX5q0rv8cLQ8liFxAxWJLZPuZWBx2UWAngD9t4IovzG4F1IltPF
SNxM0z9163Gs+5Uf9kUUWXi3Bfdsav8WG5MIuBF7btVQFMVlqLGnaJizecsETafRZfa5OgoHkKnY
xj9MiijPcCoxcaCX/9BZetqLFfJgMeSpLkDEBU4+z4yfOO394oGXHM3FcurXIvIfomzC//Vm1D1u
n63wnZiJDaQpM9NrYHlqYQIWuQw2XaQpjx1BDp8APhI7I9yndZcjcwRFht9qm8nFpbjD0i+6xnm9
ALn3HIciZY056TBmAM5QMbFwy8WMT+Mt0ibq1OI+n51kYrKDrbaYD9dvBXxldDHp/P9j/cM9xDYL
/to9f44Wh0RpNJ7TvimunpJY1ydf5xeWk7pRgr3QI6xinB33lMXxMUVbQrwn1mee9BdkvlVkPByZ
+mL+larxTBaR6kbsqVo7DOd2rTMJ9EiwLkzWMpk+3owHBmon8MjdzmrQGbAFpuH1K4yDodTQ8TFs
86jkzfQaHD9B8FzDQydiYKPyKTMA0QJoqqCcAqQ/2lMfuq4btdN33JqwudIC5GXPspOEap6PVDj6
NaZARHIBf4gaXBDXFFgYjUAU5zgSH1Pc+9OcZMN44vBfk+U323TrOLjh0X0fxLXDB5WZZrhrQZCO
QTKGXqStRu60hLL44d1tvWaMB5lhc2+w7eoclbEfOdgif2JgjtzydKnyyqQLp7MAHeosx5KAS0BF
I80fFxB+YrrExf+G7ouFx7053D8aUKGxYkWmaJThKxEdJdDMV3sXm1vsMLGMPghAMdc7qiE9g3Ss
DN90ciqOWVagqBFfN8L2BoElLErwPu6cy0Spx3wpDatPsQHeT6dBtKATS8UuZz6TkzyHhs7JpMwz
x3PbOnRGm8j1Q4cNiT7mclXTFrQUOXtxbVKZ05mxJYyldraOShAYX9x2YqTuJicqd2q38b+QjcXT
Ttda2vnVgK6CXwjdv/BMfsjokft3qYq4JYkOYj9nE6+i7vDiDjmsH/j3L2IOu0/dmRtMQnVZTXM0
NbJs87WbGwlImHArHGVhIAiUYpwOz7mrgMimmBmsMWBv0/fSuXJY6vwqRhEF24KC++i+Nxnna9sX
QAseAnfodxHs8UaK/Y4UuVdplZP51wcNtpO4NmTohBXjJERzRrVQPvjJSrpOCYF1G5VcmrPWS1R3
kTlTaYGxLIxbksmN+sPtl12vb/Ae3Wfctsts1gy1aVEEvYrBA3w7/E0KFWOBzukSgeZFan4xFM0e
JEhyqbbkv9Q9ITI90zXU/7rpV8wyCacNrQ0s3RCIFirpw+GyR+CZlNCFPp6KvwbuyAvaP/ieDt9j
2BtwozdnASwJmS523JEM+GQEJNj9+FpYNZJGDJ+Nirhe5kjZFdDQ2BTqT/11KF9n4SPhS4FCmF1H
Ib/Lwp/Hg6hfz/wrFj5de4/gtQ4NJXN7zHOZAWSeWNrNZb/L1GrWEugz+T6D3rByTRUZygGgyCrA
5DirAM5zMmpnDUez1Y6fNNzvm5LhdzpjFNVSQxirhdVUMY0TvF/xBjemdJMV3082HGJb1VH6vJTR
68E/jcIMdmS+wJw6wm3k30NIYAVaghEK5czPsUMnbXcF9b1DgZVzDNoTOCfw6jx9jqZsUE6veOAP
D6KAmgU/PJE8yLg84RDOF9zxxoKSLsma8JCjAdtRO1cLFpfA0OUmk+IdUN0ubuVyD1xfDz5t2txw
7+VcJodIb/6IftswdWLYsSHKAE3GPpn1xRI1H6nF5E652xgkzx9ZSsdjs5ub2/N/QB+BUx03QfMz
VN8NMFTt951jZncIPKgi1E2Bodt5pqXvJ0jcY5+64Rvri7ITgf1x5zIKKSwV+KwUy8EwnJuUhtKO
Q0GdJFPTdvvX8RtbBuaVi1jkmxh8sWfXFcltCwm2wsJ+vlzEvkM/2YyFoSnFuPVAob9C+8ovXJCN
jCSbJSq1ouHNh7oETtA/HWiIYERel9frRF1ASgNlsgHEf7dsqiFa5RvIjQaNuIRbMk2dGFjg10OW
6T2l1jgBHPH6Xffl5h3GUMVsnC3JO9m4hxc3/RBTT99/5aNRvyxjPj3zpLaejnYzmD8CdWqlCbqM
ImCzscdL2F+LbCotKyBWfAs99Ozd57PeDykCBol9Ft8vUj+6I6SqQEdSby0kRNtf6Wt+jgJEJkzh
AIffGOspzg/CD5pHYisZsLRdJUEsre9iZxWzPIm2HyuobsDaU1TNnKmC7mOJYk42aDfwgU6POWnQ
ffo4k5Theq9dqJG+krcUHyOAFdNUARkP9hpBJksKN2BWekrxPD8xBqF4wczzEg9MBbW7yuQC7d3K
/s1WGJ4wdsvzO9557I45cSH4oxQJ34J7XJYj2GvdYnQUMWXVXhZJnCJdsF+55PHyHJo5o9wiMV7U
f21El964p0GqEL7X7TOGi02w+Gu7bbv8nXnniu6tTb8YhUyX7kliCdA1R0r0M1lzmyTJm7AIhKZl
TWOwy8Pa94dcJ/YVmO+vwCpIoTeSpxZ/XyyD/hWJWSATz7eyyWhg5nnZOKp+BU1knQsgvilHZNnC
VXVLUqQJ/fxBVpWLKhTvy/hdLn2pY5laqjuyxv+Gixz0L78NkXbFHox0DL9FpTYcSVRBlyPoRxov
TMoiapH15HDuXCHgbz3Lg93vdi+B/rIiUQQaoMPc5E7E+9r1UDlVS1xzShk/2l38CA6FgCHH4N9q
FolsMdU2YxTuVCaqVTDSuzsTlU2F+9uYbl3n/NFAmcNfcF/vZ2ir3NmqM1z55hgiQWB8OwPl0+i/
r9OJPTk1xMOl4bPiNnSoCmVtsDrTWspbuZumaewVNNI82BdQAbQzsuYi28v3d8PtEuZad0M1wsr9
oSYaQ/V51urb+rdnczIJHZMBBuRfU4ZLg999W/znx3xvwmqOOQjvjMXxbNVjUGxNk+4a1wniQOhr
FKvqum4vZU0mRlq/EdH4uL9C4veFpdXhvgX4N/kav3e/nHWhMzELwvZRq1tEGmCBH7UBZ6Prq5QE
0QukopeFuVWxAZDcd7Q/fn8WPficTP0e2QKscHpTAcPQ2Ougi3tUfgFXe4l6wu3Cg64BH6Wwave1
Y0sXX8rUEVLL2rmA+6gibaJ6GJqsPwuOnVfSkI5ehK1xoOXOUzKs15zC1MAtkucfEW5CCIIkIbW9
nOIQ1n5jLEulKhgI5T7fRhy2tur0uXVcDDaaEeeeR+e052z5nFyHKxSA/JUfF3aC7v2lNmdMkzJj
lGbAU/WDjBG+agA3bmRsLdtRvQg4/CaqKDTjuBOe58bLmRfe/pZ9ryZa9jxyPesvNuHRh0xo2MGO
5akuXcDdd/SXTdZf8MozcSUqiGG/XKcBwEWuBIgRMJI9IAE4gNhXCwYDS4c1VlAVOUg1h5zK/pA6
WcuNm4eEkkISCUseYLdbItlUUr9sxKTPtkkYr+p66QECan/zsi6rKYiZK0L9KWrpLo8OWGHAo+N8
7WHOkf92uB38iO1MXNSFLzNGtgexKzQgaaAm5G2YPabWD0HGdmim2/poLt45g9aKip/5VO5Xm9YW
ZCI6o98dNRGfgGozTTyNvC57yD5XtyovP9B9og5SUxRFqDKAIyBpIuFPA6w2JjYKmu/mBtVUgTX/
myOon2PFGP8mkFrmjo7DBwEpATsTKE5wZ2Vj1AxStBg0xE3QS/ODBkMNQ4Y9wCrenIUaTlXl7Jaj
uqd8+sFFoyxdeM/MPls9XLiSs9GL846iPIE4S/n/0HJYcUHhDFUlrp6AXuHYHUgR6HNfNG7C5aS1
U//aVUCH0OgYh3L3P0u3WpHkBRyf+FukeZMmvc3Hqov2It0/XDeWHfo5VPmoUBoH9adVktGPXEt0
x8cgye8deq4gI3HKm73IbcqS6NSB3dfjHxh41mIlQqOzNsQ7H1HO3XGogbYOM864xBX9a5D2Je5t
JSOxRn+cgPbhJcZDApy8m+W1GhcQCZUXmwrZg7Hddim+l1ffyL3+AffcvBSU6vYRTdlENioIrf1v
k0t4EfOU5ZZjg6XBNSqqtGgfUK4qdPX3vVSr7+8FYmxq8UyDpsQamEgY+LkQ9WIbSL3tvl5LJEZf
kMc+NjL35XS8jXPcpZ/nLsEQESn0rAc9RvPNvVgNFaIXbH6kf6QSFDMn7wChsY8BmKdIsSr9Kctr
gCd8fZNZk6731dLUNJfEONR+z5QTyZ6RxOF55D70XcZMXJ4IGBb08O51EH2s2N/plUQ9ZNxkYqKf
wcTgPfmeRlxudiWIA0u5boqLJ1ggFJC/9Qtzx/mJiruAZogSdeEkKNH510nw/30HX99Z5YGbL7KJ
MT9IZNeUOSj0dzDPO0jzea7geYoAH2vtvect2PeEKgTvyuAIQzDQDhzrhtuTVkj9Y4PFmipWrYYe
kWeuFPyXH6uEjkK/rzS5C/30AnT9atEF9AKNIWjFmRbzI66PjGyV8acvNOfojVhFJxihrSD93Y8R
GvnytMlb9meuI0umfaRVrsFtfViwS+yK/YDSGwgbzSOyi226U4age5pBOOeWondHrWc3wsXAWWXK
jtpMUcEXpJdBMiajJh866gSt5Ug6CQUcWbrUi8rMjdrKeUkIjd9djaCw6h620fbvccyHbQ0eCERp
qX1wohDppOHc33S9sDE+dVGC6vPyONPpHtY7V1kso1toQ5jWorqkRKFlGYrLEtUPC/5TPMgynSUc
m1P3vzKMS4Xp8J+j2oYBGM8VvbVnwLp2ZPebtM1kgKJYwQqojljdG0O09SPMrsFni3tCilXDl5YJ
vVpZJrgBZgPdUmoaHs8mYN/e2J/i6HnRgxbTB9iUrAtxOJ93dhSzgWq2oBXSo0DKRL9iSSvSXKwi
LMfV4YCdB4B4PzjuPs9G2fQqzdoZR8isngPMdcxzww7Etm8BLoIt7ir30tX/7mS47hcT1lcGe3CK
466tpx3hhe0LkQDbME+TrMtTFjPKsWHEiqGoPbo8W9yMo+xQPWlSIltakmbJ1UWcVCbOSLwAHLSU
27euGmDoetmpbrrBLYYoc66apC4vi62xAFP6HQGoPXC7DySBC4CdnTaKriL3NHPKl2O9+RRTRUsp
BOVvyBPzuB7jh16lBjSs5exQkZ6kROLFG/S2wiegv+ZVa6Dl91zA0kcABOW3wKXsKd47tCzzEoxj
eGmR5MrEvqLQAKHmb06GIuJBMep0PkwS+Wm6sfFpMhRa3aInBYe/+8MrhSvsY5VEkVh7limFdB6r
lGUkHlXDqN+GnSnd+juByyvS+akywJhgDia66BcJl1ZBgLSzf5ff3Buu8fV6FCMoYDduU29AAdPm
kjMtbHkuAI/20HC/5JJDEQp61rINsXbkZudv0JcEUtSd1NZjadw7ASB4u8sVwcU59QClE+bEsJ0F
4W9PuDhVPW17/fj2W6rpksz6AzrOutZizT9HPeyrcXwEffmjlMa4TunqFWmIvHaPraGB6NIHRkCz
EbsreNRQpAEPXG//Ryrrb+Qf0Jmkt1f2wC7fbvAbDuE6xxwJdCd6QZM4MOKv4CshgwUZm2b8v5NO
omBnC7Vvxpc3f4gRWcev2C8EMXqQ+GpSFZ8L6HEFENalMWWOLc2EWv0w5A11E4e0ScnG3bxI43P9
3EdLN4s2lFgahU4lVXNO9zU/9nSJq6ONRgfNYZZEPjHrf8nkXZxILmpOz9X9JIUgDR0WitPoJIbC
yj1rtBpVYY6mdw/8qOIAmmihm/7NaReUlXeh01PyedrQtIWgSEYMkx6jSRLBn129aowvbQlD8hwh
p0eV2y5ZBQK4Mr4E/1NK+sd4Fq4DwsYgXaoBagXwlJQpP8dbMCNn+9JFBzbWpYFDxUvbkPgwrpaS
5knCL4DI/rSpCAkeSOzTeAE2X99bliyD8D74JONUwi+SB1W6Wb0T2CZX0v+B81KNjmpsMm8gJ/BV
3k2G1c2xIM3+/XWNSdyYV4QafDX5O0Coyz5xjL1646hjOcq0Jw0sEmyL4yxAdmnNRjnPjc6k9eeb
rVUDPD1WdIwHe26kwDDSETimF+hBcJUuG0cO4oSQ53gsOsu2KUMvCe8sDdvMkrPaJfpD/1ndTCOF
VCJZAg9KB4+DaX4N+L22JB7c+UfN3hiMR/rFsJXIRRP/uCCedNFtUJ43rxwK4HfBOUHhrvoiT65F
SUQ6o/sjoIYw3Y4PYV3YFCo9k3hjOAya7TDU0q3crHSxNedU3g6df3Cqmmc1eC7MaCmd9FYBtrZt
GXmkZAQhzrcqU41irDQGpkW1v/HUE4+UmixUCAHfMvRk5K7FW5h2rwSa0lEM6M0eXtpcpU/anrAC
yQ1m+ib1Hxa124+QhXlu7G26qQ3B+6wNFTEQprdsq094TGsgEpMxym9hRu4xCPZSsx3WJtaHzbRV
ve5P5QaKVfr4kLj98wMk4YGD6yVDj0zvtLxwl3Es3zofK6VXwUnNVq6lnFDhyR1diXRbawQm8/H4
3CQvTvLOCw/lGvSjxzdie1Kp93pQjqNMdoqzLKCdvdk5+VjupmBYDPvq8olu5WFZtRWx646f6Bmi
SPtb/HPSm8FsfmBlKENwrTKH0TcyxeKqkaBMsvQWpy9dDSxfIzb3iLfK/X+NnwfygL7FH3Vm96el
VynSt86ls4DVApqI37OzCn3akXeMPtnk0dOb3SQGV2nUAexhVaZLvWxqyc0od9FnSMdwpCX5q7sM
hhP3RPGr8jMA7ozWjNZsfAyNKWTbXEfZRcHEBMOpgCp35DG8mE6UMtodLAIeD8x5wnezgivbhQv1
TcrwyqxsPRf7s/GnL7bXHAgZ5e/htD4qgJLc1FbWkZartYH4wcUSAqhW+q6Xqq8go6lxBzyRy9yq
hOSbPRBOUfoQm9YSe2lZi4pOzCFBlTw4ATkYQ6G5FCXwV9X3Sto/wIb/ntpGVpxuDTZIg/mCDoOT
jrdW75RBTQViOQpLsnyGbVhbTowFWxrFxep5Bi6WVwIS9a0M52/bK+lue52AlAXN5i2JqBooIwKA
9dlKDCmA20e0MBm0gKCHGQoaPIbcTbgJ5tXiudYHEF9Mfj1o2Z34R/9H+z4OY1jg8iMA2MhzYXXg
C3RQ9qkdHbi1Zv/2/P5dQ9Tj2A8Q62JFceMmdp9dCyyW4AxhjSfpON8fbCIqS/uzxDMfxVRKyoZh
1fKW+W098Y7Q+3ltZbwOg71CM0dHbxZDH178OuKAG6p7NdybLbIcjgUlanHhFUCcth7+HRL0jw6Y
r5YgPuV9SvpvRrQd5BsbcmQq7nX4oi6dbcDYUH0coDHhyX4cTq1nZtqb1i3riMu8gOPPNmVmfmsb
fx9vfMVOAfja/VQ5dUYaJ/+jNqG6sTWwVAYRpVuBEfuaHWM/KPw/jVTVEIu2UraTjhjzUUSNH67K
4TaVfKfSu4dx3R2l8zB8JZWYgZ4TXJdIfsjttuBiinwMkOAqqzZO3z937Op4Bb3B4T9TpKfp+Lvz
3m8CEcA2C2NRyG9510NBTsHmne6jy+VTEQdtlOtbUDH01CNdUKXp+OjVmT7n8nyeQryAnSLfU7xC
nhLAMNBKn0ghiDLSR+94/usgriEewWB8JWhTuvdV/GvY+/osoORV7JAVIJbLYAL9NVxQhN+6kJ21
w7BvB775pT7Zn+CNq9rvQk1yId1/hRFfRhqi8RrR0Mk0DLOkXW6vkHwHdbvqoy52U9NcxAVQjZON
XC2pMHYBp/QTTD1RBYOu7B939jKWr1R8LcceyvmElFavLvRsHbNpTVqjQ5rP4c9NOp7qD6mXgr/2
ffYnxY7QI658QJZ9lLGHbkS/1Epz8/2sW1koCFkzZx/BS98oNv3dCAj7ExS4NBv7Af0nhF6tmdNd
zVDCkATL6NP68URPF6YMSYpn2LfdjPqlSB210cbHzznwROVNoLef5ctdaH7+i7c88xxDzvjU6sUa
lqfXO+nstFLwY4aPv1lA/TAEODek+ovQVE+pxl3l+r0OIVWhqVPogxJX/wmHJ/5ZuFJtpu5Bv6TS
SKBVlsY6QHTRkrc7AfKEn4AYjFmMXAYTB75xfbxredpIT4gy+ddMp+KY3ZxpIt+IcVXLbPnoSZ3y
2/mIOyong408OFmoh4pDHQeQvDvJGCzA13BhgEhP8HV9dGRMaA4DepLZuXSBGX5g9jXpTZIfbqgk
m63YisVF0ilhUaxKwx1m3hfvleCY+cg8ZaTp+kKF0/QAVor20DEoANTSYpU4aS7XZPcs6ZXHTSHK
jNW9KRwRhsIa1SkwZzNRAC0OdJeOaS9qx6G3OpHKw9cytSOHio6Y4gUIDfPqrtVHc95XYvGzJQ3+
vnbuDcjBr6CyooY9+xx9AApbd7PovpYaswwwvpfjeUyY//tjATn1haevQPdXZw3UxYx4jaPKjZWf
+JU5Gxw5GPPMfMk6umPlu75+H3fnIKFMYsukkhC/hRerAmUp3vzp+l+SRKvyVO6p9tSl//1WT7Uw
ypu8eTutfobLLDnwfBc53CtxQFTCdHfvtlUR6zXI8oTvY5EQfdSLnbp4Tk0K4omhWH3L6y2ktOhE
cMQvVbYsWDd26hd61k6pcErRDYHlUskvs1O47DBJ8SwSImzJSY0pVOQokn0EfqDTZfdXBw/0KO0j
7AnJJC4RRsLl7n+B+aPuK0RRrwIHHOcmxr2KqF6kvOEY5s5yiiPR43zI425kargm5wucnOEBhBB2
/kts5QRDeFs/KP9zdGUsrOqe78ORsLir9L2vGHrNh3lNWLyMVtXIqLtxFlFcXRegkpukf5rP8vn2
WWt3iL9YJQNOk8JaKffT5gGhfZHQS/NsG203F9mWmxY84X6POs+YebNWIdpFBQsLAQe6dOoMSKqK
Mq3dkqZ+Yb/bwXxy+tf1upjkI2Ro68SgqXKScdK0gt7KYyOC+L3G0H7xvqFa3Eo4/zRBVg5gb8PB
AYcz4GgrHHLuVXNPab1auzGPTXsNYHm2P6zmP7z9Jzhzmn8GZsxL9/tkgPM1VAx3geHigjQO7uO1
ryZKXns6EwYn+/PLrmzPCOenOwFURr9akPTmU/EecQ54k1Ut5na50abyTc4O8OBjqg5tyv3FRpbF
tdsogjoq2aQmeav/gwT9wrvxzL2JXQY4XaoRaCXmxu6bJflxW8KWxhuLgZerhJin/g1GBPss5VE2
1J2KBfyrqzNzUPdYFsFE/UNCXDL3bI30TQI0IgXHXdoxQv2KSEfJ3xKcdVlWMUlceFueSsuNA61l
I6ganxJIFuF2XX4ZnSjCa0LoKpxiDEx+KjM7gzAKLwskh3XTwOj8At4FFoGfO2leZGl3U6wc873G
oe+jQbm940BB8S4l8A0ro2ipppPDsGax0J/NdiYfHhxLmA6EiaE7n0/EoqEqDKpJI3BCI2UluVGn
dO/9LkJY75PHL5P+WA2D6sbdfS+hkb0n7Bz8n9Lxv/fDtWDcmZdLkgZaOG3yL2eeVWsVr9gmnfRn
TFzyop4xP60SvVJqKeNScThmbqDARWu2S+Ztrm2fwuN8k0UkCy4W0E9o7hks8SM6u+v++o/xJmgG
tSrAEBH/5FT/f6DnXLrAV1Odb64ndQG8uFqUs693kF6OVmh+C5QDQa3j1sezBdBqCcYS8545hxN6
TgBDyezeUFJiXcjOxPdsfgyPKgGfyS/2WkWsVDmwzhgvE43EDaEd98Ijjs8DCTQLSLYJdOwkfXL2
B/8Se/nImAwNSVCWefLiYrcV/l8o134e9ypeomFJPjRKBo1bd2Csdkd0Gjgf3HfcvtoI0qcIfykj
mi5zcZico/1xINplhmJLzqLGpKDzmOT10QvWFd+H7f90lnuq4kXe9f6CwaDGzqza7c8ZaDqTxE3c
87b7Nfqyad9v65biniGHFiYMAJisvN7RRmSNQUKBWJDxlgXsDfSLZhzdJc1lSUf68OZlhQdmQOIE
UZT4AcVcoLthW7vAxI6FyAIXyZ6XS8DsUlVxITIR2NhrxrLX4C/2K/HnXyioorwKDHSB7qoUGqGT
uuRY7nj7+uhl05tkr3sFs1iezABtDKRLSDVVKGAg46qIllBQ6lRKRV0v5y/MKb7ccwTnDMUoLKkZ
Sdni4W6whJayEpwAsqc/cQ4MwK4RAAqO32AcgUtgMB765xQSnZ5FmB7Cfrg4JUVv4h7e4+yrNdmL
Nj598ernUbAVQNww1JAM9cVz3Pq5oLTEWRiQVAOGq5bNCvsYeqQHkGmf/g7uUH1rQxi0TP/fa5hZ
UYgRksjyPtikV2alhjI8FfhQmbKpUvK/GsDORj5vUJBT9L2KvIzzlz8w/4XhEruRHQQgpRGdxl2Z
CnarCVrvQvVar5l9GTMVHXFYF65m/V4FqF0GkT8lFTxx7pkPLL7niwl7LfZqNUpyZs0luPNqT32e
UdjeQFHvZgg1yfSiwrME3t7EcftxRvz52QznuJqvp2Adgb1Yh8fcmP82rxHxmWObTNZJmL6TBSj3
t6mDcaoeFsSlpqyVTCgInsZLCamwD3Ei0UyGVERwqLbcdfzPi3AasCVf2MMYbmTfAlRMJEaNHUYz
nhCwCMNAh9aABAQZNMPC/WDfbSu4/QgiJjatXLaIKvJ6G2w5MBcfTl+tUiqG5KGMaKpdPpoEp97g
m7dEbWaHqpqHLFCBqNW8cyrqkZ10lx/2V9lRslsCNNPzBrEpKft4BJtakFFJG1PP1l169VsqgWJw
gGH2EW3Y8G9qLiC27gvzYXzGCktIe0dXFlOvQYBLM90o8fVsH4LUGY7ifL99/5vHGDjXZHEqcywY
FNR84QNRYjg4kmlFyNrXgm1i8qCBnLgmzGZcHl/7e8a0SpYd9bL8jdO/ym3a1DI6naqI6gZ6ZmvA
k3PQf2zY9FJNeeme7C8IJrvWJCBMsQ5IJz4zLWBXxgADevAmBUJSMmV8eHMistJIVKAHpuXP1nnU
7h3pzm8j9DlNVW8UXvhb/I58X8GReb6AZD5+MDWDvob/uP11mRzbOHGpgMwmWFOPzwTutNDBqNTa
2glsmV/RdSCkE1coDUVbZPvo2NT2BrW82VrTZ00YFtzHyNFV3pUoanMNTblTFAKl6hLdDnbwuVG5
T4N06hnLN1UZvNsnNTqK4pU/G6MFS8J88aMMBYUpIJaQnPS4epXDWIE+XZBLh1Pn0UIneR2efCe7
EVnCnkl6DCX4bxlPubYi4U0PVTHOEg5zi7GEJZk/5Kwq5bFuDQTQ1Acn4pfMwL3lL2Dub6uOxUPt
GJ28mR/1kJBDvv1SOYSP9P2l2d5/gC2/yqOEvo/w3EI5cMFZM5z1NjIv65eXD+mifkWkKiIxy2kR
qteIxeBhy7ncN1ayguOD0VYZWHiMPkzTauN6R5N2Am57omsaPvme4B9XheGCZmwtdWtlcW1wY3QO
NhcHqsHI4pBV3xx6lkrIXrI7IiVudejsbjNlLCxtyyLBtAMikMFeOr8I+u6HdbJyAIQiEQebpqhS
26lybX6FebRLRxuQ3JWFMrfh4STzWFjGptxDXnVeL1yo/8vUfh4mb8ik8dnqHtOdXKhvISbHYuxB
Zrye+GoBj66qc8KSvr8MvukRFW8dd/SFD+8h6+g36URpC3huLJUdH1lFLyqgEWhGpC+RlKPXMSUs
CO4VZVVqY7hKijCxhGdi7JevTySBAnOZhBuUR8lCAKMFc1hDI+Uq/2xW5WLNpjfBtHk6X3iM0Sf0
KJRnGBgjjht8XQwQF3uF+JjCLOVxjRyxVn/LTSpJSkn0HBcHwIG/lNrjWqyYmkTa1GbZMV2iI0cL
3CPWs3I1uBdOHKN8cQSdNA0ExCILMK4X4H9Vm5692jLLyuSGf4HZne35u7L4gExAxFYoes1/yU2w
3D7sv1/X7BRjYIe6PfJKGeYplxSHNLB8FSlhxj6XNvr/O/CBWn/0/Lfqck8ZC2kWjcQTWDsTKAKr
IIqFSlRkmaBQYC4s8vIHcVneT59blqmshH31JOr9zm8QJKJC4pIRIy0Q1ACbf6svR28UdJQWlUsC
8w5eJ/YRZ+ooqGj96+hdZHhTG/sTFB3PApsTt/+pvAbffn1WX40Bs49bQXV9/vSnoHj6B4HaaPsq
O6PsRiwVsvQtTgUZv4bsMdrZFrMwPMloPp5Ree+HVpuw1rN97v7FnoMCXqP65HVFyAmazQPvPq1P
Y8Kba3qI8eKWI0TciyekOTFJZp6EwVV3jCuAxmV3IwOZlYwPrcyW8LYYXW+WFmvKCOenD3i/GeAY
ZDDlISVXm/Jr4iqssyUvZyZD5qNhUTBZQ/sVK7/c3gHEOzgLaP3GJ6Y9OKoZXYRPjXhGKjd/sCKO
pZS2CFURcXWOQMmWgntBCqUNZ1lmOva7qLdhS9AQVR8L8Up3i9SAr7yRvuACY1e7/D8Z7rNntQ0l
7BagexJpQh9GnhcteJNcwrYlDbyrEkWlEtFyR5yWgM0QajP5BKo3/slE53yPK4cdBnz6gNZb2hZD
2A6PRg9EdBPwc5gJfFQZ1QhuLVAbEogteHNSTYo/21T3EfgRrl6oCRxsV/OSkVY5J9g/RhUYC7VJ
Rb1nCPb1l4MYxt+oCwWF4zM7LUeHEOOzrZcRUfI3i7XJFvNA4dhDffGmqg0Z8g3BkjXWJ9WvU/Hw
bCMVp1RNPLFTz16/JE2spr6Xyw9JQ+zECchcryceOTpH6xZL8gkrt6b9aTzA4RQM146ibc/KZ4qG
v0px7BjVwxhHFuZsQuTeKGxDQIIZQkYA7K06hUEZpjc1WoPWxDIkSlwlrfzZrL8+HFHqGeLnqFBI
GNlJM1yFEXk0vkdF71lrnGaTqkPvzqzIFg5L3BuwBWBG9f1VlucX/fleWiXwpHBTd0McRKgMY0+p
nzfgHF6j4/ZSIw78dsS4gBVFrfNUgNgROGeSlxkyEJT9dssB0neRXHLKC7jvEhGNZx6UF4y3rGdj
LgQYLBejKgozGo3RhVPI4UhPN6W/NaojDrdIkKUQ0C4GRt5Ja8mI3FIljNtke2QBlMJn6n03QUKp
uZxCJPMGwkTNND2TGqcPM1YTSlrRwZETQIcFgqxa2JLHRujFIH+HQtdqT2fKfbVTvTnzPI3NaTrU
2OEEgXv+FYDzGpsNi32lo6e4JO4TPXgmlwUWs63ZjQCO/XY/wTrqEzKGJRCiSqREPfkH0BzgSCsI
gwYQtZImyCrLQyEH8glzMb8KSIrGqgy8BjmQtEC5qIdYJ7WAtEFDqvGQSkz9Ax8Aa86DO/8sR4fb
EKC50GHUXpHwp/QDjsLP/i9lGC3PQy3qsIIPNVTdczbWWwLgZizibAIDmRoN7bpJrxzZnNh9y9mN
6bSakztbB3JDMO1A46Xvg7kgSbhL581WM5S6wsGjRaKtfPNkegYfaXctoScLqbIZRM2Y0Wvq1oTs
u0gkk41IWmMsPsOl4z3i49/fk2w9zcB27v+2Uu/5132FPWGgWzMHuFyekuHt38s1limZUCurDWmA
/zKa6B8n/NavBn3LE9RMeXJgTx1IryNBUso7Uk+py1SKOthDP7bvXO8iHvBlB1jmEPPkUSUhgPtq
ph7qCjH/5oYftcSZCJ1ZFYaOQxjg+eSqISsMucObTqn6orXtZ4S9t9JdYp1rGxufg/BqWF9nyV8y
lna6IZclrSvMv+Etj03wtNhikRuxEvfQ29qGSbPAFrKURQUAwsRqRxDx7sh4bINOf1VOCI1U//Ze
YF16Io1YGUcRIXsUzsQvPgKrOws3KM4gp+pnzD1sg8ib5nCjye3NJ4oUoaIRX/b3ulcFfhCvhLUb
DK89faz93SOEe1F1G61tt2MHI5o6XiM2VXNGej/7FIX1qGpdPd1KsBM26fRVEjxDLzYxfaN/tTQc
FiUGUmw8NWR0NzPEvJmvKZZV5v6pKJ/hcOD5m171heWCgOmiRztWh8fAgdWVCJwIl5b5pomozCMv
ore6sqQWaZo6swJW+L7071mKr3ozv0GsaCr2eObjbN+tSYqg7eippuBTgtl7Y3eCRZT+AXHatxg4
nz1M+lgXB4TdC3aGM55KLhSvIwmMEbtHNUj3kN41gMpKt5N2HlNJZ8ef9YqPz2tYxsL9CcqEIGd2
nMRRKB9sTJek84McTMuuSTyt5gLElO5O9iql3y5PRED98CZuElYRGxrylZX1GOKhHpYh2rvMimXt
1iHRuYdpgahpy+UWefiwtmPVe134kBk43qC2yFibtU//UrdF4aThEa3DKTGdzucLCJpylo15SjFn
zdm7gfOK8EGdtebeeDbPRj06PPTAptnfoCmd38UjvxEKHzeWYmob6t0QYP06Nkch5hILLmIXUZXJ
6U18eMFUYNy8qhPvqeTRNFn2+UqQolf79ZrpuwsXqpGHju0W+h1UfWmerPxj9eOvwcsNtQU9iG9H
sfrXz6ci81YsZkz2zsCXBv0UKgNXF8X88TnaKHHLxdLgB9WpXCefVd8H8bpCtaknYP5HaYz55tcb
7f5gPgmDItjn28O1ndZGLEmTEDD5V6nedYxEoCpV2LgUOV7OSjP8+83biEuz2yCQZrhDVUikrsUw
u8sqIr3rtIyAd+1c+dR2Br33Du/olOAHCFHs6eh+fR9XJtbLwUD91w5/H0pH2NO9LKRZaqogKFV6
QxEH+M7qJAJ/v/dCNWdFTD5ZG+W1TRSARSNuoqzWRPjGIa21XhSngHLAXYHlOFlTFJx5RSOzBIne
jOftyk6QCNh7KB2HhuXE5qD97h9Fg4OUSGnK39IPoR8ok1TqAZIp2DWnPMnoKIPMfq6lSmSmiSss
XkPEEs3ydCjOlXRD/czPB+R78RPSc8IjPwAGitT7N1z/AsvCp4lTWmP52ygCBnQzTL1otRknm9ia
XsR3l+evI34mjpRcHAQY6MXsUfcEfon+dNLbMh32nIluefjBoolVvfOnI9bh+0dH6t6nfr5gNZGI
c74S+LCxz+YCJuuGc7VzVnREgMw2deU6KPczHbJU0ruO9LboGzyi6c0wfD4G2UWgcNBUYP7PHVid
ixiXkOrVJUGGmFmGv8jYiizTeUKzVekwB2TwhhfaSG/kEkCFw4OUbAwrm1Vzh4dQS67jKLQtvEtg
k+JHhbnH31aN0iDbo+O7ThhkNpaqLN08lhiuB3l6wL4QsBYRvjdsZjlqiZ5MERuCI+0rAyvzTrAU
j7Jw6TQRqVli97uRMA7OBjHQwHWRaoOMsdq+q5NBPFe9lnQAYYE80y79id7SDrrGNuUKquwbGKPC
/4lN1i/rPoA+A67LLHHC4GgUbHlzx6km25wyFHvobazSr8k++d47HwiQ8zIxaadbdHXuIo+G/9K3
VSqxf859SvXxmZh6zkhNSXsSCeA8/YIMdZ+vNte5bh4jILQ+EBbXWrVFwppBD9GoTcv6zSpZa1EJ
WdfL0T+I/+/UYH/Vml6ebFcMQvJ23wSQaqvK5rlfoZO8oXKG4Sr+66YwgqP9tmKL5jm7Zz0PyKjo
k18qXk7/zY/a+zVRl9L5M+dFaeH1qMNEB+HE/UDbHDFTCtjd+XNAAYMcZP8oycMf4pWGXUXbvcLZ
pNGR1oYXU32N0Ui4I+2klCf89iLeNeBQROneqYPJ8TcauaPlFGFnhIXMsdXTdkGpbMfrwjD8ECA5
g1fLifyG8eeFmGAyDiQH7UrlFqWA/kEw8TACRcnlqJofn85772rV819iEGUDYKenWUkbrlSZM/dx
OEesOpt4t/SaABoGrOwwF/EfFsD8x7HW/LWQ+KLSvt+DmLKpRyY1CMqkmi1oU1hqC8sDZJ84cDzp
OS6724NqmaA3QZ9nU4VzjEgRLBJ5foQsm2fzfDK79umREs4dnWnHdK0FLgR9pfv6/AYjQrILr9L0
K4v6bnJXRDSdYVUPkYXVZgh8AA7BdXDqMYvMokz8ZY/6waz31PQfiW3Hhl6a+bUjhBagBNOBTPEa
iVscGVuD6dfqNEJyKK8rf9AJrjUJhxeEAIIMSn3L0TeFWxcqm3o0Ntf/po/92PaDwxmrtDnWV08N
rpxDXKwrQWHcMYN76i6wSL7t1k/aMPYxEz5i9qPjvU1Jqbk2XwUc4g57VR+iJ9dz7LL9QrjDv4Tu
/D8CvzibNGHxJkrN/Hd0AReuazjMi5tJF7EwBa6EiLCHZJra9GbgGPNrmeL7hEHVs5WuyI8Ss2jJ
LpadN1eX4pvDAg1g4F/PHhMOwMAZ/FNajJ8hBkRT1W/EydsISzq3nTpextRhlwkKrRwtvethNg5q
Xjo1QTFPMh1feL974NqfiZ5bc9r6wIyhzQZlOKXem1HIacgwZkSZdHWQfWBuskqvAaBxKfDKBQhh
2DHmJer1V1dguPIfY0W0kV1H8AX7ElhuPJWFqTT9kl1cPeaAAD2nPS2fSk02vWdRZU4fwXadOSd0
atGQZeoEfTm8d4gWLo6xtLSSar+LuuRC5kjk14PvifkiEvX5O4YnoXQhuRnCGTXrG1GqDdILXc5p
SfgqPrWQ4fN32UEjdgmudMdiqZlhUsLR0YdSkANVSNVw1xevzGQ6OQr3xvtfsiheDdKKv4rHawaZ
Dm3MIa9Dznz2LCmHROQBoxDrFWXHV1V9TDA70UHBnsjTYaGEC5jIqkJNbhRXDCSN4futvjqLWbr4
PiKRzuswvntHF5ct7hArXDE6NrCUEZuCJzmvl+vtfaIiuYSmjjrONVPBogPAdOBKk2ySQvZqac/i
OCoj8n9HaG820bH0k8Gb+GVgow3DR89IXbN5bH6E9qOBQiqYBHDaRyRpBiNnFDO+Vs+m4KOzSovi
9zyfBz9+Snl6IjkNtUX21OeFwoZphExj4Gfpg1uPQ5GMsFstjzT9Iph5fvRgcZi7uc5zjaZ+hXQK
q+7bip+31kRypD+X/xab6riABJyNpV4z2WNznaYr/GUxnI9oBhYlzX7uhzXIMEF3W2yvPNG19/zb
dpyK8Syrct+icfj8jagrF+sBkdbnS7R+yhQmplmxt0IHt5u959tU3l+xV8W+JX5EBvDcOhtUhYL/
L++z04aXLblqDwA0ubPYTG5m1gsrI2WVY2MWXx+SA/UZ8CohdYDo5xGqgTFw5wTN89OOaEUPD0bF
0R+XXgRd1M5OIS4LrZK/rUp8AguT2I91nEJNC1d9+QZ+mFB48CI9lHNklTu01STbkqD3f++3vcBO
K7AO67OXLh7YDzxmO11PNWEE6DRPWOD5FbJBSO79/r3XWz49MHkaB6nAg6Go8TbOrFt1m8bVHdMU
nn/cRSQMcOtwPat13Waam8tzmcr2V5PEpE3evyY2LRJ4fRxdst344eN8Yau/8OFlctEFIbdFzNjq
W9VFFMjnjFfFpM8X4/93dly0ilz82ZoQuumWvyxVuy+eNRWw3gNWCSbQ+BnnZqEDy94bbQ5U77Le
CcEBi7+U5pPBDBhTiUrvakjXr/ZeJbga3I8x/tAMnhkrPX1hyGsir1jrz+bvc7ODv++9RJz823Ja
ojSlg2RkoMgAxBvNP4vNQGR6Lq5w9LrwXL3GfFHV0iToIqAEvZTkeCG964MmIMBFGLja8aZIAARf
deh9Wabyv2gTPDba4YlpFmFBShoiEc9mWdQN7VeTut1xVK68SIbwt5TQfgbqA3JBoA5HLCUdh5SR
eDklWYHa5GWW423NWSk4zf8dAcI1pkpY9mXaPz+dGmkP7sSVf7s21w48iNRPDA+CaAtcOlfcKcYQ
i6VZSba6E+1ILNslt7yKWBSwj5+kuDW8PiR4qCF5zK1zHiyRAPRswPZR6qkn0SWTBcRiOpHItvXC
dpiITzCBJjAIQwZhPyBozVrMea7+iqfh/7jDzUFolZ3MetVkpakHgDsGApzImKITUEOZz24GEtMP
vemaL2pcim+SydH7mIRj1tGBhXkAc3USZTWlc2dSo8Z6NUJa2sfRZUUlOd3ZVMdrU4YkzDW2xe+9
Hw657SXs+5Iv9LXMjZWQlhdaK01NdIc1IKOKCb/fED/BYkZS2xmVov0n+Sz4pD7R04LEUK4mwVS3
OwOWEH9chLwBtLtmlL41O7L7LOsXJYj42s+X/qzTiD+mWc4ieZkx07+K+rkSBy3nsLSVX0020kPL
5gHchFG4cMwZ3halSdPHOtQnnfV/NIVVitSxsKfFr0bEYExUyDBY4uYpCVu5KIB45/i7chBq9bGx
IGn7nPthfSvJtyZ+FfkoCRrU0djbby15FM6Y0tMDgE2+Xo1YmEHuMUxG0ctWfK8N4vWM0Im4++Bw
yfs9Xu3Dxy8j1uV+Gvdc7VrxTAddviw8HnbExqhPdMZOk2RQ86t5Wg2OHUWQbdAiXiu4SAT4I1Kq
Gwp9ZheVIA+X0IY1X2F++vkIPoUR6CE/txNIDs2vo93zhv1zQfSQi3oFtmG8pIxWafcmb9VU2yYb
UnPcpe62i36EuuM7gs7X2+/ceYga5m9xN7p49jk3kV7PUkw0tMhDA425RGdkzBy8RQkWBgr77y/U
iBu/ZLFRHUie5D20YXPb5s+2+oRFOYOyypC7M8I++V8BjXBpLJIF0wBT5pg0HVmJTkPVy2ozDm43
inXmkCTaXEJFy9FVxzxe2aCUNVgiAmU/yngvaLZVUq1L3S6udRK2ZwpUg++F9KoVUSY4oVoxpWDS
Af1wB8BwWBXjkfzuaXfH5kFJ5rxQLMugefBdbOs+VNWq/mZ59WjctTN5yILfoC4102c349I+vzVW
+CUjeLg0ysN28SxmaVm20OQlRo+A4MMzPYFvsU0tflgnVh9/Ou9H/dTCWX2yWvJmkC0EmjUUXVS3
9B+LtU0mvks8V69xEyrhAlk3yyHbZPeiGZTsM1krU38cC8nvBlve3MXnXzJjbGIdNwko/5txrxoU
EG8yoDwbYAdbqXzc5eEEQMJ83SEg/L15xjkamMTUgWAkExIs9r86iLlHgP6xoLp78tjiMqKUOVTR
MThCqVapfWbisv2MrhUDohkpg6n8MlOxOo3Xma+ngs+kMzGIkf1lSwNPn2efKrCHlA9oj0Y49aUo
ybBaM5fEzzyrgrtuNCRwoXA94mFLpJbscJmZ7ZxnoZfuUB8bBTUxHOPolmI+cO49AeWMMGb4I3sg
n1gyl+VR/T9mLASPPKBsl887qwnrSFBqu3gfzEbiutmVMWRcHLrpvPBQC7NWhn30lCaBjUBn5gvX
gSJtidTQQBlr9HmrJ9QadRH3q1mpaGFV/ruQYhKdX599A+5dwl5LAN1YZrTTrbAR9eh5GBeYb6mB
fDUdJCg832j6o6MNEOqnGtazC2/zsZlV2HrluMNDkiYLyiiBsSec3Cgo8XqGKlR+jQHnnXihguAi
u4lsy34qFkr0oEtrsg51wVxXyt2uEUNgPTJvFr2t/QwyDYPea8OE2721JsPtstK4MVZP+/LW0JIj
bxAtpWssOk8IyEK5JnG0TRYhg7D2BXOPxwU7pX9JVKOcWZkHgGTK1dFy1HwPLouzjfc8ou46xAow
7/Tr63u42HZ1ymBC5Mbuq8kHOytqtzqKu6n/b8Ow4rzigPCfsmV7E7M8VFAxBGz8fLZjsGpdjSWK
5zaFHcFawLdkVSJGsi+3hgpyVvWK18HQt9tvwgYUAymsZgLTb62C0NYGO3uAnawi13rQTh28OxG+
q/lbY6YH0YT2jqZZnRPUFj50u+7hig72m/LkAk48M6ywPTn+lfspxU4IPeb2G4ObmS/RzfRax9NV
HySk8+ToI3+FIHu0oAoynEQhpfJ1FIAwyBv8UwGAnOiUouEbQxtpQuBaz02FpSsv0hUfXcq1QqNL
8++dlvOn96FPt7mTbDWgIUAvsbkDtWnlhnLoXgJdBqNESUNTL/DknkYybiUUfWey+sYzhV3vTo+1
Qm1vi3q1ehGTHL4z6z8s0ygbgJMXfOVPRAQZ+WuSexftyTb5gAOILyTYYJyswNLJqbXOofVNJkb+
FpfvsnVwGk1rL/rbcZQ9mJmMgtxZeb/F6YxKLWAdPbZsHSfp2A4EfZW+NFiNVEQY4hNZwNlCiSv/
qTWspLyDUiBQMaPfwWA21VKXcJcjjQ0SPsgI5BFNzhaWyV8PeSxqFlGzLRWDWxXfe0j0zDfOMVQD
55+DZ5I4ppidpx3tUj4hBxtiMshw0H9PSIB7KfW/uKwGSsdOFA0ydluKZLch9uDRKntJ7t0Gzvab
fJ9328jroxpc+ae/gSsI/smIHK7BpsxVLBvdFN1cTbMiqH5ajOFRVomR0i8cf13nr1nYZD819Rvg
cyPcRTG46yEyI4rSfOmOb1Phks25ffRRtR5UehpfU2inWQEcKcTBpcwSjn7Ba+e70sdtNP/Mlnhm
0+6t+N4MirmcqzBjyAni3NiDsU/KC3oXqSgyxS+SGE9J8utxKQi0GlV/eM6xtCS9HC2EtMjPalLz
HLZqn09ehuq04Wmn1iT0wSbDz4g6g4EIqB7UzNLK2tGYUsoqoXkMo25i6hswbR464pHc9mcAhCl1
YM+o/TFeXhpmjBZgfRsRkPIDbtdeybzlgkvvXxYoUu+4iD86xdc69+Z1rJf9/qfmaVx+EqWeJzlL
P7B2E+pFY4UhRyTngyOdJRQyxgT45XG9pzmZ4sfvTmmK8gGTb4Mkbur6CXfvE2qtFiM2yr/xUrdz
dZovo2cZDCL8RQvnpRyxCqUs6bsKmVBSMYL8yjds2OAOI2Ut2HfrTNEBUYR2tGbnNwiWQpcupdb7
ek6wiXCylWcqigJITROA4OKUfEyvO+PE9nl/qRT1NiNeMPOqFdRUl+YtYhzCrWZeccqtWsTpTtJR
5xYVKp7L7H6bJHiyymSwZYH7MGhJ44yYzerJig6tI4kTLTt3qG3J8LAHNj1vw+t4653V23L3mzre
IZAQm9Q585kIFQdNhSnGGvPv1scZyvorUbH1hM578xtPwj9z/MI22L95XCT58gW8R5K4DiFcTdqK
dyuYPcVhYIscVdyrw28vSkq+BAEFPrqN31QmiMDwlknN8WeYhF3rqgUgYs/A8WGoEovhOIj/EDbZ
nIehFOIyO/yG9d9zStBhQSe8zlJefaIDh7FLoJJCcQ58OSgoxeIPkgQtt9b8X+kacVcskqJZua1X
v2D+fSe96v8zxgsIZV9TQmIZNG5lPU82zogN9BfrHZFVmvsgLcpUDdjSf5eCoQ0YC7oz4GUxlmdt
vB+ZJONJDuAHvKpLy61ev/PIvQCvYegFB3FIto6optxVWQzljFIVGpRE5/xjsyKAJb69Aix1+6UB
uLJ5wwMQPVEvPsp2qYJiTc/vYLe/WJWzpSwq2xU6KkXhZfvktUbAD4GxnfpozEJfIDgoXx26J3/a
5N6L5IbOvcwSevwz7mRDhUg++ljjr+ioJZKUnGh+lrCdS6heyvT5RLysK1rRkVoPtrAxXr7eKDgu
O6tyAO6ZGhSUR0V2Relc/X/bpMEKL9WDGdSq8/QGFjkfH+7X5FhGbGpXB20hhF7ooPdgAlwpEy/w
9s2aCp1zBjoXe4Mb+cykILByayB38EPA34/49TMcuY9hTg1PoVRQq77i/GISiOMqWy7rgndH6afL
uxEhuY9TTBrZKsGQ6G36LCdBtWDEQC8hocBvFrigtD5MRWZqtqItli2Wmpxc26GHESvukeripdA+
F0ObjL3QZ5ifJBaQDrBXwuzWhKDySbVcBS9bQyvW6H+21iAGjxG/IKhSQxoZibhXJ7xcpMXKV4BW
MOAtBKu1ueYXvBK4TCU+xu7PU0acGcwd3S6tbmtyelbRJ7ruPmGOYHZilI6XmuaF2vaV5qf2xo9g
7KmVoUs4Zh8i8hl0kOGSRg31tJdHqvAwuwQcA/yshwBQ7benhfqsR0zR9KNDtD3Q3T4JSyMuw/xj
ZC2V/lBzZQT65Vx2AqCSyrwda+YBob8UdIZzGH5TxsOP7b4eq7qgM+ZHFF2pR++6hjxhwLJ7bQ3S
ZhydnKYKffBYVU7R8GG5mYMUa8ejI+6rCN1DNHgP1sNtiC7oy7WhhGBH9FZLGymXHx8BvnQHCEFs
KjsD3toczRWxWpY/cZmOrKxSr3AHeCrR/+nCbCPBxQ9HW0wDNpQ4Q96CnMMzyUrCCdbtq4CX2bkj
SGOIbXM8lf2ElNAPOQFYKmQ2EHbMLSsvmK6kceRtTLHNorssbQY+PnPN7MY0Y44z3CzWkCVRq6b/
nE+kWSR2L30xv5kem/9cpKZxVvJi+F3cSyzNQzzx7izgDwGcVrkk7WEY3ypvY51iR8IVtmjbF2ZG
R603GetyleD39SvR/ubepb58GgD8+j0yN+6B/JAKu6O0AetQpWNJXN7MDcxDKZTVt7nlXgyEXsK5
rE8NjBWPoZnIBAFcW5FBlisesyaykaB0ZM2ADwMWsGBRVp4uonRuXtoXNDrm0JTTMo9/5EW6iKTn
lvfeMLG1xNNTwiCi2lncT5wVpTGFPhIIR7FyNydCOxSOdtqM5aXkcpkD8+2urdUj3vj+MODrlQhr
QNfHtkzZ92kHaHMRnoKKWvzpyXoSJhqHgONhQ44HaAQ62URMff2JAENv6Es0eFYjst9y3HyH1tUP
I4HboirRCWTZiSQTxBVcfpF1jbMlgYzEeev+cW6+rTZ4QAZPVAW6kv4Kn6JOBZyISEVLLs7Wx9l0
UodN8HWi1iCdS1TdKYoWtnrTpit5RpLATc2pwxzSox1dyuwtluv5lAem+g1tJ2lXXvfzIS8JzvMF
yaDbBAbf/0OEHKH0oYrN7VzjbDf4KnVrT/SMBVPvAXF4o7NretBFMw04GNfrBUgOwzW81jhGmfWm
f/sw3qfcI7+N8fzM0s5DvASlnKEJmWMtiqTW9PhrxGoNBSW4X4mDaBTX1G9A0jcZxS58aD06IJth
M0ZVeGmWryVdepI/CgMFbA8m7odCsYgMYbNKn9d8SH8XFzlrM5AUo1T7wu/5YjFLZIxHvjeKP8Aw
0JH6IcyIcEIemQ+zRFNoCTjBahn8miJdWdU5MvOv/wlDdhE9CGmrepLgbI2iLggYSZWmlLiw/dJK
N5xe7IItKtXdtePMGaAHyAWPQ//24kj2buqnvo1bOpLQ8fASUeAlfeeIBgJ66a3kRbLdnD7+oi7p
tOYsH6jh2dEAO8zAB6qa4RjTWzyWIbM86/ppMIS8l6eK6m7C5iugsCRbuEyAir5eFOXoUNZ3Y7yc
BkxCuI1MQIOM0JCuN74hKNoqN4Jsxlr2lnmrVnYES2t+oc6GSAbHkVEtMQyed8gPfXlpcuiLwQuO
0DeB1JsLj2nhY06/cG2F39gj8k5vUg9Ohji8WS0jfnpNDkfMxBa7lQ/2e/26xX9fEuRissVr33Ca
6WPVP1IJpQgVjz28Ze300kaO22pr7a3F+4uyM8mNA4sjmH9C6VVlKKGHCwqOR0l7FU0S5i82cXAZ
KDyqmQ/0fe3ok755CoAhKIqubrnPRj6z3uEtUxre61eueId9QUunPnkQbRgwcB/yW9c6aa+Hg5nl
uA7i8xbZTo5wZkKm743iHOaADMlsQ75ANpZOo1YLZaIejb0415ldwpPkyk64x2hGwcIYNs2XAeKe
+PcwERp0S4hbK+d8tRigcMS5VEKW+eTOUzHgOjaFe7zyOdnk3jkbLwl5L3dkjuX+rL3uytU+SoYR
1mhV3TpmWYTnZHoICJt9UhFHxtZMhnyEyR6BrSGakLW5nILybmhrSgLBANaZXHeGrxKzvEXO8Qn7
fZcZkXdyqByv+M08vyXNRmS6lnRYq+fJNpacx7Trr2c8SV/eXc+8b6Mt0mzqOHJmNcUrayPtt/QJ
aVE/HaXzhM19xf3cGHfZdQTbpVhy7ZeFhaAkb+5tsHrlAK2RqUqimQPRSR0xCpN9x/Jw4iFZ8k55
oyllwGGf2ylQsIISnzHT37NVegKGdDNLs6t2d/Skh4/8Ie/4w0N800XlcVl5fKTdICh2FHtZPxuk
QEXzsY9tR04oqZeJ6jSVwhv1sZLT78NMVPJy+WRriw4BDNlp184F8cQl3+60k9JzQemv3GSxjTxl
Hzh9QQATeA3ZNjWbFlXSdiwzgStkPPY5E7qP9ucQJiiNl/xvILU91TKi8Y3MhFJCP1AU/c8BoFCx
n7K5FHLYRFVq6WHMudv2AeFLXauFIITSNisl62bzN974+0n10yaWF0X/DEuMEndCrPUmSDvvT4wc
Yu+HmMdGrGMzBvBNUSj4jBe52LuVy3VL4mXPZpQtgc74cCGYaj/uY5ff50lsKwPGNp8UA0JbOzsn
lcPZvRxt+xPOPdi1VteIsUrFyR7DbmQBbztRmh4cxXNfMpyrUltioCLfs+FIl7lQUvmxmTVYmUs0
vxsj8MfmwEfVJ7OBx+QgvM0C9/ZLN9CU1EgYhKgtMJUTeugSnQjXP/Y6P6U1+5M7WAKfldXuJ9rh
nsBaGATVx2fgLIIn222R9MhUz5Qruxo+C7doVb+pMTleEYYEPJXua84ChGN3osi7UVAXJV/0w6Ix
GV3jl1i1MxUe3u+CsV3SpFDxI3Pp6al9MfrQeXMY5PoZGjxfsZIWu6rCmoTUvA+OKptxdmGutkco
KqJObuBuqSpbN37mXCO3Isc00NQPZ9i2vfZyn0qej/xnIMViNFAnNs4yGpSM+z3pEbuXfAukMkZ7
OJ2byvj/a6EWt7jmrXIeNEzDlEzm7wRxTu1i4IY2fsxM1/B2QKoGkoZeNiLsRTnorWcJso+StalR
oincwgeuO+olxBV7qTvAydfsr1PpH2jTI3K3flPTmnr8gJeHeyqD0uzqDpSuJzZuerD7zLngcAo+
c7CJjDYK5WCr1cXMCmFAbjqvUT9g9Cf24XdUfiRK2cRd7hMGTT5Tw0QS7h/34ImZAcvE/1RQt6MH
PDkVpvSn26mWmn/u+TJztFJSDBCajQGBF6CkW62HX0flda91wKxWdYn0S7xT8nSbDKX8u1ICZsjN
3VysCdEEN2nN+ebD9/u9NaCfDSv7ajzW6qD6TeHYvVPKg1KsQz1zyWftHN/SKhIBFk1iaPLmwAZ2
p8Qf98Snbzm3vdLgpLURNNgiOoc/8AGF1bkoHCZfuVG5H8B0jYTLenP97pCf8CBHH0iexodqiwNG
vqA4FNrCHC3lNnIvf7xJakTusdxeGWaNGfUQVYr+SWBSzFPhh28h8C70t51KsPbmANxxPZK1yQKK
OhXJSc9d5ja571Lybq6vf0PSEstJpmJn1sjrLDb3C+kyNkN8hkCqskkf5Q0tK7La9ADnXNsMzteh
pLp616KYkmrjQArwUQLNvydKqRS1EvXCqzDDQDG6ApMtPFJ8OqDYIDnB3NBTOX6cgRqmg2SCRQnx
Maoxm9tL3oS/DfoWiKeQpOYki9y2xQ5U8Sya7O1aywnFSmOjYtOHy6CWaK8+cr2cxw2KUz6W8EHW
cZyWNQI82F8gh8023s8F1W+ZnHIL4ETojf7D3sHTWbsd/zVuIP6KSsoCbAkdy6DWLquCTVpAy423
tVZ20vxTgpkywKDaJbv3hYLJsvIYo5E2bv9R2Nh7FAhsAB9qxKB+VBIlqrnFCTUZJewPeV5oyCv8
JQesLS6hL7Izcca1QQY3PJMt9t4cSLl/BKo7TXWvJrzy8Q2NeLEGncZQ8b1yI3E8kAStCWcDanXa
LnYFQ7tO9EuNHpt/CAssyUxtGss8jbkH6kBz3e7Y3SqBkFNErlDcUmTQ80iPMUK4RQLsANJ79C4E
ZL8s6B9CaZYFT9395QCcY7bhMQn+3XKOJhp2qTaStu6fZOrdYVTgOkezq/I0A7djKFkFI03fc/XG
GjwB6FTenMYD2s5l3+vmF0l0PHv2vDFLK43PWup09lklnZYgkH4KeEXs4I5FcJTMA/rtNFygxxfL
4r6i1yc0i0Th9/Mb7lcirS/PXqA6zV5mMlcKm5MtZ8eEv+WYBoAhnVxVGrNPFly4yMYAvCvWlSNU
8ePnNnNwpB2DIEov9R/LbRkCWkjVml5PCiN+pDH/FAxi+Uy8fFhf1QrYR7nB7tfhKG3qgXrri+x+
uQpEUJWqDrwWsnxeYplAhD5Cs/CuMS55cXKE0OGUP9iJZkmT41RCVlQ3epVlHo2McyREASIROHre
o7OLTL78zjLD+TAr7ZnJc8563Dzh0EZRVFr4QHMDxYnGrg+VSsnJxt1BTZ5/X8B0bs2fIDcyeV+d
zIY5rLSz7NOcg4WXih9zF1mrsFifKsbi1WrMuJdoLZPHFZ2BtUOKrR4bep0T7tw05CqdclZczZ9A
VTmgyp5wMtGjbpUcRYRdXHYJUW7T/xpGULwGuQr8fnJMANQJkleOLipOmd+cuasGAx7pfUFhf3mj
X3IBV3vPYKfottDpbKnIGVjT380xhR/uRnpwZdoOCURUK/XCL7uSmGQPHWDHj23AmW2h6cgj1PbW
I96BMHkTKx/NpmOsmiII8EI/F1T8js0HntaA4SfYEOppkL1CGz908xQkajP7OP02FACjbWS+N6Hn
A9O71lCX5tJFpRB+HBhSfkxYQDwVj+3oNawlhDsfUHdteWDqRSog8ILpHl2GOHrrNs9b8AYraQ1a
IEdzXnRJPrP2eeZO9X2qavLn1l2RzwH0hERKV9nQpCpN+1vhqCqvPglE43IJi+zr/jIpsmSZkLJF
FJuNvIy4YCTj1FxWTKj0ZOhOurcYCs+Q6kFfSkZ6+ruxo9XOjzLwBgG+5XpZ16hrjKYKD6suP8/o
OEEgZTV+wN1tkGK7Nzndx9E4YDVc6Zd2LX61BWaP7ZWObZrQuZVdwuUfPyMKijv4AXFQMo765M0T
HrbVVF159m26SNn6ZhfSP4cfFGmP6X36fT9QNa12eQKJJDzBDhh5b4dHuzQ2rP3yTdEk2+deOX1K
Qt/0/n0FbnJ0X3Lo7/0XMIbHxfC/U9tsAd62DJb2PaQDPXN+zuTpFPwZv0ZKdg1dKCjqCaMeIg2X
t59jXZgercDyaoMa3Uyf66aAmTo30UitiZdgH5NliUrRZxCa+dtDI4N4FvrgYqMOKW2JibOPEKKW
6vgx5Jc/np6I5IIUDFtEOYRc/KKbDQWMLbN9XUquXqL/9aBezDW0+ZbKSQggibmA4O5jpGhCR+QR
NGegtG+KI2AYD1rJF19C0KgDq+fV13XXUz9wYXDHi+2NbR/3tBKynRmZn1gCug0XwRoK6D6UHaRn
zW2fEQVUh7RofF/JSMuuOHDELmtcMyBstylfimiK2FNv8FYMt/fK57stjES+sDEBMU3IVbLZCHZW
NplAZAG/JlkXWi4MHPQBtfHh1dFdhhVYcYi69BNw5XC7utSYDJrl64CUOeXmS2pw3/ElZWu9sm+M
TkPacYOgZLF1sm1Q6EhObOaxLrMtmMqbk74GwumdYS04qD86yi1BwmjsuofHHw9ngJwSFZVWWXO9
8mAEgmxBWPs02kPstX7gRw5NW7OtcDi/CMYSphNJEbRYi74lmvU70up/5pvAPiKUlQiJcBCY4DUV
ci07/D6k6ATu+lpHFbaWanO8/B7bH/3ypVmUrQBPAEwxI8B8xwallIC4Q2XylyHIQMpveKQMqgId
TCNCVngfQDXJWCq51Bq42qHOnEWuUa7PA9jsejZczz2jYLSeJx51XPamfa9YdjG/8sY7CrumRLv/
rCXwSHGJ7iqdEFF0o1BSpRWz4mP0YLX6kA7712STk9eq5F8FWpMHowUKFEv0EsHOKj8n+3SRslZK
GMt+uzatL6ICusCztqxXWVlAcfOLQWn0x1adHfpOz/zMKI0VxzSEa9p+M/VtzL+oswk1To36wpdl
zsHwymjSmfmNLApLYzoAfnO7Un+Mobb/KXB1R6/pwDVrExeoL0i99v+cQ+LhSQQiPaDuz/eS7Mgj
uueOQFBKvP8BS7rU6jl7U6e48ZLfmPiKEs2Y/PbHmZuivTAWWP9twxHLoob0URtMpfwNXoJA9Rxa
nXc4/wZ+syJiedXQw0dIf8GbpukWrgpqEeL701HHeHOSRcIv8Ldp60fQnGh2NfXGdqOYDjEu52b0
6aJR7Wcen59SxEPLFUhhJVmvG01bSASXXtyY0DvyzHOzLLgQKztsYYktr+PoQmargRpiQ67jYTrP
ZMx56UyF8KCRPMN01cOrZg9Qhpc8Ki0mm5BJJdLWnaJhnvr7Cwi827kUDZ0wxXiMd2UCpLtEoBKT
vnrDGT6X9qgBkbpsvS2202J752bW7e+/WZ0G/nyT2nA2Td6xJJdwvgWoM9ccwDNLsLfFE89ivg7M
Gi13P/EvyTZChzfs5wg+2m0Ek4q/njRSIf4be7kLqrI4M9O05ZomxxB3zRb/o4kdkETDqheJen8H
mfD6hxt4T0jYi+4SNIMQaDEuJARt2pamN8OJ6je/GdxyG3m1Hwef/1Y1CKmJMWRR5gARtJKe4KHS
/iNIUhMNVGJAW6l7Hz6xxojMcEOsSk9G+EHFM/X+FCdEV0bMKU3e31O9FOchwb0sg4/gHxqMfHd7
alyr5vzxQaAcCNNo5cl/wrQ8HOJlXRe79daFCOgzeR9uEiDxb/nHRZ85vLZtEo/Jzv1/HsmoLNVN
9VzPUaQAb0vWkD2x9L8y2aTYElS0C8k/OF4/uMfqVwvKIlRJXKeJ7EV06JGaG1Ulrg6oCqC0BiFt
KZYmafSNPEF+L3v2DSA2m7HXsqUF2SJLvzCmQrWcmHfbBDe2s0IuDmSCfju+0ibdQGaRwtEy7qPa
dqyHHcs5fxjTXeh4LLoge0IlbNEV+Vl0hfbR20478L0hvZEXjomgEPl8YDABqeE70TeA9Q8f3yXU
TBt7Hpgq/CblenyJgTwjhCh6XT0P3W323iqecP3krWrWp98IVqU1+Mtu1yIgaJwtEwtAyxNFpNx2
KCE7SOgZh10w1wHTx0j5Q7WBLD2TkhZjPcVJ2Mamad4wGg7DU9RqvvthlBF6PzfrwfAfE5sXzHQU
6Et5qSBFY9/CGJdJQTTVAJJ6Eu0/HlhskhFBpFFkjcL827KqcUQ373ADgO+fBuAq4AZPhKJsoRPF
6+ZZyWzhGM0GKmrtt0L9Mm/XlsgsXwSK4U7Ub8vsJNpNiF2vp/LkjUIwHO44HRJNcrOS70Xftcgt
FcNaoqQAUBOMfVANBODR+cFcUsfPf+lkkn98S0oOtaM4CvtceJiYc2rEvFI43bQg54hM61BX1+6h
5Y/pbPSS037D4peviyMNFM3vW4POps+1CF9ohihItYVkaUVf249NDSeO7XpW95EPxsdCYvmQF4fG
V6UYr/nURPJkEzQIJ6kBYSiMDhdCOQMnUQ7XxQNiPMhBuU3QsGi1hIiMxZVeCh9VUMHsSr+/p3Yy
ZSmkJ0VyN8akuPrFwnDccJKaNd6NYzzmlokQaAE4BsFSWo+0U9rIPIhDWkfLfb2hyiu56ZJ36J+q
P+MHm1xd2iTwZFWa19HP38HjIcAEm6INYQHGJnGqE+Cp5QK3ofWAFBFcohz2I0saKuuiyfq1RqyB
0aVgj7HrsEAo8gKha2/Ckf5OvmzxLxZ2TOSrwKcIaBJORbxblpTIg/l6qlfrnzVlebI9wqM0+GN+
J2//w4SeDYYINXNWYGFQqoX4GGcW2b5PLnnbwibmsYpIc900SNR7P4G98g/IyTWJrI9L6Pybuz5U
k05RPCKjxldmsk5RvZFfWOWtbph3qUqGaRt2Iqf4TVAtvD9ALRm+/Mey3gBnsgqXRdQg0DPwFn2P
PmJMwCV6ZBZMfzwMch9ql+TAG7uRiWXg9u7IbRIBmOYARcBN7p/arcvVivA3cOefcy523lYaN9ks
xCNm6tkXdd/lfB9zMNc5nlhp6iau0R3pI9c7B8CD8SfaLG+vPxsFxe3HEAbOLPsBkRotJMOvd7cc
MQrylXscc3W+MEUhWoeNv8mLmFD4+QsYf62LWkjWpvG6SwhCkIE+SBAQcfQeffL+MN0Ji71O0+zV
i9xk+h5LvAdj2MOc/NVpyaEaghCIkE53VWPxJQqsLY2DQ5SjBVjfFUup3DkWJnTELpN+32bKCpAg
lOwYV+98FLFEzaJPJZ7VMOBplL9tdFKYQKT5OrFhSG9yA7WV3TTqNPgp+HpBrZgpWhlVeUO1LRnh
4upGiZVrHiIrhaoNmMaSS7HZq0Pq3NNaUJHjUYkoACMWokP3/SOTTLgKszgjvMMoo5Aa4Rd1bten
hXaPTnYByzrCJWVunrGpgJ5AdJ3SQzFqlNU9TJ3LoeC7mG39la74t6KLRh9mIExNSQ4cdJopNwdt
sOrj3RAlDh1SbBTxB/LPblnbA4aaGe8oUgfMuvu09M42R9qwJdXz1pNnTbohObbtf0nwMFPjM6hI
ZzbN62RWDXgEXozUx/ezD1zqq+wyAfWKX3UJBs2pWuNJHXBvHFwdTyBzp7nLPP1l7lvtTXB+YWDv
BENsRqNqU1oX6n+7kFsKSJSL6MgG+24EPbzgR2JmSlYBa/o5UtJN0ZN0SLWv/7ubc7iUWS0RNHU7
nGIj2keFIBrgDnHYbP1OKzxjww7spDoTPey9AeO6OhmRRAScqct1d2IU8Bce27gN6tCedpt2alEo
Bbs1Mwn3Zz0GkUKFMSfbDuPuPHyEKjDhPKC+OYjvPuwoy7dQlyAMg9RoAqmmQZ8F+xckyZOEe6Gb
cc/ue/avD6M5hq5toULm6m148xJio9CjoY5bjjWJmHaJmNTWoFs/ZBh7K2dMOrS4cKRrweGwOfqd
g6cueYiFbkzMPRhDLSmBjUEWvw2SUAiycbM/8W11DwJ2UXEYBMEYYK8NpAHdQ3b/31HDLbbrpHmp
zix/4Hhm0clou1vc+yM6fRdmUf30q5ATkUIs8XoOKYAPxXsIzurju/jgb5cfi2Zy1iH/9PS8UJr9
kvbGODyTaDTcddiTxxfYKixrtFyuqJ7uc2jOBJ05RtC8V8B120sm49+6m5poEvjUKU/YruKeHjUw
xuJS3ZVOJCGkh68V+wcC6wKCyb3Dkjiu3uMheep79OdwxMfFVFI+uS2BqNL+SD9g4g3rrpT8fRff
928osnfC+Jok9GEim96uuI0YTu0Jd4hNClElRwTwMbK8fLNTVqecF11Pfcu73ymyuTUvq4D17F/p
EKNqfxr0FBQFJYmH3AFkjJadk2oTzp9H6f3LRnEdj+xBkTdUUq8VN2lXKXkvI/BfhSg72TUPRCS3
EVobK4lLBUJe6UTjP3tJnzxQL5LvKgC/HFMQgbWTKy/kezxpmsmCCJnPnzh6i8QYFsuLFgmZxE3/
gvALnu7D86w3fdgvYM4adbo3v8mLPrlVOZFu7eRdl0zJByHGG80PvHbtnlpO0QopfGgh2jR8dBta
3dvxTMADCjV0rAArB40SZxZczZmqKHmYzzomAubHbzTz2yn8Ta4fswEUYKsjoCEuGTrNpBNTbycL
jI6tFHHPkKBKLQqpQ5OoMSnLSZReBFMfisfqJ2xtJSZ70sgKY3+QBYjG9yYbR5+skI7WX/LkCKB2
kvF4FV7U5URtklOUb8+5owW/H4jRmr9/K2d02scwmF3HQDg3og1WvNJc5VvE4QmfZha5a88lZTql
BA2/GL6IYootcRr/Z3fAqIlJYF+BiHCewgJ1s4LspII5CkpHGPJaV58D9YqeS+KvopDZoR2eeoO5
i+SZo0CjU/npIH7mUPV5ufL78LR6/uqdPNa2zdrxRon2auoiOapM4o3bXq9zbiHBDtQHiuvIjBof
gd8oNFvn74SWuvWu+7fHQOV1OYMXz0QR6weVDGH1+ClM6kmOz9A0eFg/I5Vib3foVK4FdfFpkbk6
9ShOwl6G2pfC47Gud0FbfF7eSHFhv6Q6EydJ230RsMm34ftRpYNH0NNYzv68SjBl7AZpCCbuMGtM
Zn1wRnNC3pcKpv/9VBqEtHcmEi/cRu5fAAjUlzN3ITTA5QsPT3PNB+Y9eC+LTLeibXGeKvuycqD8
ZLeebbCvueSXFq3T3fDI2QhJUeKTkO4/L62SDjQRC07jQazPrapH98uSJLutT+UT0419lfJScECc
W0bh4X+Q9PGca6kB98Aw9y4ZY/ej7i/cnACtketYkSfLhLKiHBiSaUJj1atI8oIwDvNLFpg42D1W
pzWknvhUElUkdBaBSs3Qjd+q40JRG8aviUA6g6mZSHLN81KqsttDw/m2jYAfGes0ivT0Fq7XujqW
LBG/PyjiDa3d0U4lcccIcRQHe1ZXmb/Gb+5w6RiRsC15BbXmjuOWX064ONOLwHa58832/tH0uayK
qk91Sd3ovcSjpPvumJ5oviJW7eSmYLGtNy/hus4IzS3cZAfM3DB4wX++Z/RF+nEiTLk1ZyAmI+iu
L7pEJtICjuiz8tt9rAHe+Ho1/QW/d+6p6R/IGVlMxGB8cE29YHJS+enmwzvhkikTv85dOq0pWrYC
g2Lrdk10HeQD/Igj26mpWBrjo5I56xhEI/wAYORuBY2tLdynHbwX9CntCPwkE4k2DS5oCpnZhJbC
c/gzlQh9SONiOyxi54DYLW7SQWsfjYj3BBWReL+0+iT4KgjT6B/+R2eohuzeo+s+/VGJrV5gkejx
UXCbNE3Sw/5YMbSBchaL8d33QsISPSEYTVEovDN4vJuS6gPkpvg79w7sKDLRtAXysfz5EC6D2hgG
AlYt0Dpd6G053TQrzn/jZBa73xcTsqdB1J7+zdVHQklK2VqwPL+xVTDA/J21m7Rm5iafs5Im9+Ae
yhLAJ65odlacr20BAw7Q/59m8kLPGElxrZ/Ud8tX2J1ds6pLVPx/9s5v0mXOFpxHKI7c5e06c9K/
0ZrfWLmK9TicA5i8eBRwNDBLHHZ1oiCs52zLJUD3jNwSt9rH3VKMBqkYbDvKtSjsdvkgi/xlbsE2
NgdqXlNHhoRbt2ApIKxJuERi8VS3NUmKDQCxcEhFmY4gyeq+Er8rOpdq0ftqMVqPb36PfUgxyVBi
VIsLduyeBmu7YDNDgl4bMKlIdKFbvQUgIb7BvkSvpPVEF+HG+h6eyAbtpEZwvZn+BnxON5IPB3Qd
y8EL94Z4M3eZk53Ng3ZYU7VFtJ3H4B9wpnNhAIiPlgIvpy/gCwes2dCNdKPesnjdsvRlGqeCtp6k
h9OCC6AeUMlodjYEkq9ivZBV3kYiuiWIoqO85aC9Dy11S4haeCXuCQUKMNUQs9rsqL5ProGFfP4V
qeQ3H45/yCPBIp59hd9Y7SJ3jr3DFnJhOeY3nBqcWRkz8W9PVwoIWsQvmU8mIlhuNSwRYEPzu/VV
9HZLsMDCgZgqKaG4lcqFtj3MaAT/W0u/7rIIdH+2Q0Ki1EoRZmA0kdY+VMJgfDDr/ckhTlGjRS+E
m4/w5l0DOQLCRG5GwTU1/SBrqggzc+Vwpp+xTBCEds+uDsUi+sLdF2e0VFJ58yKcaKxyys1DedRB
zykkW+9pRvGoaVyX73mK2o+1kKnXs50ZYJEHVRN+XsTrDBhXSWROt0HipOMbwPgfOPppKCJ5hmc7
2UYplYzWod2arSWSVC2WKx1Wt3H94vKfH1FcxvCGurO5hWdd/owzqnIzAHn4XUFhfXvMficsiYhM
smmtyeIM4K1Xu+EHAa9EI+VL5hCeBvh5rD+KTeqfFvvSMImHTPySMQmTIyQHmHsJiG+9n9fFHaSa
WarpQMVMibLQtkvBQIT0fccLyviqAjrHu3RTel5d1Cy4c6iXxruKtKrYOkvBCXHxncMc/IiVzc3w
zaP7qeXFmVrwTBhP2/JHOzHilT/9uoGcSUtTS+UGbkI6TdLpijuoJyDkQ2dA4tSaRCnvew3dAbPU
8AuKOQ0+I0Bt73l+S7haUClG/WKbtj6yEEy+3HgFvav6a25mPvIETh7LZgPu022z6eZ+iZb39FN4
ZF+KIqOUyzxJF39HRjWro7H0PrMbGe+1UxfV2JrF6aJ9W8NruEkfRXaxPGWiIsR5MQrtacagdoKc
mG49I94nxv8L7XkBcEt/dcZ7b3N/CnlbTpXgIgsGPVqxbMFL6+FyqgLKVXFGQAfznV4iSMpeo+EL
1RG5V1oV2tF1aWzzLWFAbSsSXDlBeDfegglxTc9pGFxmLuwyBzT4LVcNDkRRLVk3KtA2kQo7vDtz
uaDQlb457FrKrWFDPnd69p1WWyK4jzsad1QzqJSjQRLWFbKyLe3+5iuyN2XVsYZwzVLj1Ds77lbb
71WG+sGYrtNI14zb/5iMFLF/0f3Q5Uw9W+jRBlqVHYBNHF73ky0zy8iEMGI2KWdYzW0Ygpp89Zav
C83saoLG8cFEhVduA6+hYCOu/lzFU6C3RMPxJI6VhgerlZhuZhVmBjLW7WCx4PvFumwKWJelBjGh
/WIMOc45z81rIq52Tjsp0yoGgxu4RsFlS43hsfgUoqz8acYE8cOOjAiP4+RjgxF+DoAmVb0rHavd
bQLho0yfArdjxbuH1A0fr6sCz/nnH8bQC/GQD8jxuodo9h8UQiYICyhf/mQzjx96zuugWj9/p5uG
TvaesZLoKKXcEkZ+6j7Fvs0iVPulFIEi58vWSqvgpcyAwqThrXUsYg4UFczvqQml7bRN0+7XyT9E
8otRswMe2oMaBOzsVEoYV6KTI42JBoSsvhTIgrxsY1/F3xP8uqH36Ndm0AAMnMjjQhrZIn7Z0jH+
8r+6liUzj51sOYbkIQSyepMtx/BKh99jh7c3eUoKberY3KffoazI/N4e50nc7Q8D6U+o1PJnbUie
4lSbSHaKUWBNcYj+0HYm5Y7qnbj7U/8kAEPMSzLnMKgKuMOlw3yl6VBCE433Emgrz9P1Y1CXEumC
LD4ZJ0jgtylfQd8nCuRsCrSnWEBA6Dpr3v/IslKgJeJCrDKcmrUA8JAfdcdZdjxMbeqtcMUYtOLW
3pKLt07m/MosObsjJshZKg/m0CvPK7j4LdsASrpYkoMf4DG2sdE55ai9QWu0fcSRheys6gMPpP6t
UB27WuoX1TmWsHIXkIHEl4yS/Xvdq+0NfmZmtKB2mRd4jTxTwR41g7Favti2aJw6vcEAJo0vnX5e
47NdmGuaInhKlRYRILNuEbyXaU1aYYaJiOwFnFc+f5mM12yAQ6Qr++X+2c9IRDsywW3of4oxdu9/
wMW/bbDdorvaLgY3IUhbNcWmOHFbsIoJ5PeCdNqqkixuy8dSJlqTbj+NPPM/mjnL38aAdl2Rb7qP
brV2qpzRtLrZCBKm9PjUQlgRpcG3n7ap3N9NlmE8dxOjF5EKpKVYYj2z3GzQf99zfDBxLXYJPqyp
DknRq7NAX4iQPGLc5TR2bfxGc/hKTSdDj7T924WztVYiHKsLKbhkRnEBHF/sPUaCiphDJUNVB95P
vCLHU8Oc/t+vzLQGcqchgb2KA0IVlJNFtkrpf8cilKgrxew3dfrryWhGXr7Eqq+a68XmAXzIgWbW
ngAUvf7cw0qnuO8YUT01HA3nZsx1vkxNlXQvf43LYc7CoVq64uk/6uod/919CYkFx2hAi6otMN1y
AmCkpmITtQOFQnTzGshj7qwH5HKMak0Zp55DfdZyZvq2UWdE9eMMR4WTdJ3aklKQu5oCDaK2YOs9
2u1Uq4QcUfuaj+xtXtPPJlR7B5QV1QXNj7AEtSPcwFrMq+LvTOf39+BIMRM2WTK9a3zvp7S1qnv0
ggRq7tOhj9sgQoHw/5Coy9im8c0aM9x4PD2MPdsRXJPfToksnsl1cP9RY8rppcUxHtt0dIW2rZdI
mGAolXvUlLyJG135e35nxn62fFjN2d32BSiF7VrwosVaIQqNU3ev3Jvx5SrfySkXQlpU25Obn+3v
QkksAkLS12udYvBmaNay9+ODzqXPHwAQjnIKqPWPss3sk+B5T+Db/1DBcKJSXbfKtrbUPfgLxWef
7fs1u/paoEqrD6dGHSQC7Q40ypOZr3Ry3Fj1a0eUH4ASSjyc2oJwYEekm/w1+uEHQPDyO6vihuHY
WsHgwXcQg53LvwpErKvbVUF/XtBkBq17A3wckjpx/n+ICgivzyrSs4jANrKfuWwBuXGHD/M5ZBxG
jC8hMwSh/jjzA/NqeVqJsj0NCMXDmVNZ480nEvKJkfl/kNgAHb8L/VyEkh5p5MstE/HtZ8rIR+wy
snVZfKKQRXvNdTSZAEYPYOcYUvtmjJWRczzR5v6IhPLUoeupopP8eucFGaAR1DQVTVSHXd8oqblg
wedP3X6SGdDiHh5KzUBHb86rb0BRFWpyuRD4vvJ5RCwshh6tG1Csc8UJXV7NP17Oyo1ksHl5ulwJ
3tOYahybH6hVy8pjziS9H5aMbd4hFdh9Jlc+d9gkPhK0kHobRG42WfM6FT/8PX33IlZ7eXQW764q
0y6Ia4jXC6ISx6dImq5D1LFG9m5SUNm5hxUze/y+QPKV+e4CM2HJMpPLVS2WyPzaSvMPHud5aNSj
wXLbwUBnmnNrcVD81pgJs+jT7ThW2wyfy1bgRNv0Q9ScACITXNTwiC72KtkX0+Et7EPoeH3rZMYc
2U3GWtwg5J7TqHURjvJJaqJ+iAWqXPLaubO+5wy+XnBC6NZFXN4iNipe75EmMeMdmCMekHLi3Mgc
dTJSY/YrDtk49gW3G9cu5E89a91329PymN10HzkPe11rg+kPYZWt7hQAsFfOW8NxXz1bAj/n0EDQ
vu2t21SWiX9aXtlE31Cg+C7t2WohvkKWDgWmm6YA1VUdJktcW9kT2CgUknh0xeH6MwzSq6IuJcXs
xx6v7VxkMeN+Cglvp09mFIYwMIP6LsW3+gfLhv9Cm6Y7Pxi/mPsnCZPoRPal2DMBLmAFXCUfEqOw
lJ8sNbHaNNAU1xAgwHZhQwJBtsZFjDDqyZwfN988eWCI/vp4h7SOCyKRd2KTCRQ12sky11Z/E2e1
VsQLaMSsgDlKOQmDM6mMEe+Lv0TJJKSoAJ3t03dCtDB/rVDRrUM8UQVjmx4E4rdgOtHbyr38g0Oy
sQqljSMAfN7cdcekNOpB4JDy539Rn94btr7V1ahhWaq0EE96Tqw3QYkXE0SCeevZSBtLGck/pHkL
xYrQ2QfVN47tr7dkklI+JUhvgcBcglnLhLK+h62wO0+VyOrNtTeP/Tr3nqiCLEAVkjMeTIMWWcF1
FX7M8//g6P4prOlOHR3c/2AblKcofDuC00aqur88pD7XdAEgynF37HtYbUmYDf5zqYnFFF0WxjxJ
0HdNRMWnFJR+xkFCv15zreeMsCnbA1lfiEezzKvmwaud2jUGe4y2LuW/QHCHSwfbmuxe6TWd2mdw
z4o7T026MZdfrq2GW9LJkGYoV8PHPjuLXdfLDXQ87urUZLqOXpx2Nm1CrGteiCekJtzAGCVgnypW
CNRq2+kFRc51DjTvliposDwigGXTSl4G+FTuT8ufa8CzT+UICRpYL49ipzKpMbGAbhXE7EfDrp2F
DBcJednFDIyP2N7M/VnIHC26GNcCWYUMi56uB+BsP9L+kwbo9Xclfz1jpX/s8qWnHh4g4GeTLWT8
CdmvJnvDwFxGKG4lcChF70yhdmnigGDzzejPRegvo/fiklm2xG7biJ5d77SlFCwrGSCQPzOkv3zL
KFkKFKfRd8C4rOy623bY/uJYHvd021QJdojwl84R3OVeU/YPqnvlG+SyBOmheC+bteIWaE6nxJtB
35V+JMo3xmWoFGsZ4nFjGHVC1Rnkh/aJ0zCphp/2qEv9dBdb73TDPST3qmSZRzFuiTu13RK+LZoG
xL+jRBSGRtadnhKenxdlUndPT3f33VfcO/OFGS+y5zFqyKvP6sFbLVJBpwBINJY/ewZHWzLqHaRZ
1iA5hFpqsIvUr/3/Ug4780aKqfct9QApF84VqvVkKKMdugGjBLM5MGUAj8hHzdkXJR6xp6kcVOE5
Q/fyqlt26yKaaCP4Rzy8rwVbAJxOZgAsVgjCDJLs50vWm1SzG8fo56AQitI5CySoKLygxhWf2cZX
+GzegSlWZCtCsyl9+hNUXqhHFNKQp1wPK6Wt7Z6O6thX87fPzC5WqQolDG4OdSfGekz7HxE+mxWI
XqVVT5FgzJIYAgShUZPxh8b8eIU1SBFJIAnbxkc3Xc5J+EAEJ4Pp14K+BjGqzAHpb+p/cyRgUx5R
YRT0pDAw58N8MP3qAudBD5GQm9x4EwyuTVMJMzy2RYqUb2Qq8GVjmgqEqUAaf+Ua+Ax0AVQwLWr7
PGriMw5PfL0vaypYU491lyfdP2QavBIKKlzskKh07UiNaKq6eSV+LUrLRylU6dn2cb9nICgTv1QS
WdvAnNjJCL3h6n2xCxSzaonc40dcn1KA+NiMvFIGGLfFBKlfVW0NZb8RbKOjkBX8Wx4c5XgNx/qo
XiYkEv/a5zhZ+AFp9hSig0fMsn48iPSmeXDaXXatAEcQM0fSm7+s3hVmt3ox0Wm3zsFD+CX5yaxv
sT4MLkBcOos95XA7Fxv/38wRt6XacIgmafAkF+b6UjtM7OeMF7BcKVCsgbq6Or/NpF80pYaWLtcr
dlrSaa/pEhaoCs9td5OEei2HqMRH2oFPJ8HQBa2Y9Ey3Z23SwU1fdCzGQs2I5y6ZpZiuK9PEHGOf
aKCq4+y+Q2CyLRx2GV8qmMr/EKnHp0fmRAjRLjXfTUWFasrHdz+3GM1VSZeFiZ09ymuUwvs49w1O
9YZrqcOYuvhRDWqPR+/x7DDXvLlG9WLW7oZiJPsYb7hJhT7zapiSB/YlHknFMUDDeadGG2A90wJP
/cW3MQOq42y5cktkSpotUaLYYTsVtTflPxQeOgOIBauQxVF+a9EOySBgRxvQxqVfyjW4RuNONW9q
YWXqA7knILE9h5m+T4wyH7UqkwlflgW3Ra6ehG0p6KdGA/Wt29dDFkJqqAteZzQqJaNaGXq2Dihq
dCmV+65ZHECAmcmM5bsYbp0nBc/8WoSm2mBW6mJs9Vttx87Si0cj8iCQA+4RZjJUdiNuU4O8JPh/
vtrs1NnjqAjXpx5tathDCQKa4AGK0oNbTAF5Hu+239kBJ1jpOlKAx+miHqLiQidgvam7QfBfwggQ
9GclsMZYLSvU2kqlTknrK1iKAMzqHn7XhG+jpxgf92Om52K28RzHHFNc2+7fQnW4JnB1VUq/LiGq
/j761hjI6HzOMvf9ClxGbWGxqyoindzQ0f3cwklDBkhbG23ybIFmB/Cx8kX93v/HISeSiqpCjGcQ
bWeZvhaBAcDKrEKWER30fDTMdFtk5/acv3iw2k8F+eQPdLDC/qE/B//1I8hokWnT/9FyE7DBsS9w
IPOeRT7NjVHRBkByiX62FGvXpHTDFLxMc/XW9VSZNYNBpjskUpyZE4gJf8cfqaoUQWBa7XxfwFYA
dvQnmmVyzvcmWn+iIn46fYmICox+jC0B7XXtOcLs7FV78lYRQoLZzS7BFDIIzVPH2Pl/GZqz0SsE
KPJYZ3TE5iD9mnOGWeAun3JYBMemCRu0X6qPoWOyKX86f/dtoh81xVtqqfOd2LJeSEgUmOotaiaH
vMRWEedButMQgv09fkhGLmhKNrfi74woYMypT+TZLPhNLaFrXvF7iq8vcTfH3gzjAtXuwKUpxYS3
7+ztJXiptwMBO/dcQRwMrMzSO230k5z1vbrAfwOeXXpoqlvlEJOI5y4WB757s71qjsxiXvcRYLOD
KOQsUyzTvMc/Lr6mZHaCsh5NcS8nj4qmi9OJlRcJNJilfAukEq1LZAuSniCw/tlovsAiSzbxQMJj
E3FH1YiwZX8Vyd23fjN2spP8X6ZMhPGVeear8MI7Yxb24VUwwfFfaa9CvD3aGUux96ATFsFWD+Lc
80B4QzVuKT6ey7sMRchnG/bjlGCdaHbmDdwhg7SFPCSqk0U1DBxmyE60RbpPqV8e5xieUto3cs8E
6j+5GARFDgnE45yLVROUq2g9x6VZcmEDdyqpj+jX1ZsSJt7DiPykpIb9Ra17e/c/vTDhmCMPb86z
M5SFKQ98XkvEMLtoNCFTdpTLgDT50q6fbsa9lGnbdrJx/CVHhbLq67XbAxqypmjaZAXdG4DNcKZq
KLkRO3doY013AdxbDQhREOYC3c1kM7+nlyKYk8ZXOnQ8XGEpiwXKiC14Erk8AcG7caRGRaEbr697
dNj7heUU2i+q/enHlbyzk5fgUU+yVsTqE6/T2eeaivxgDTssoOcQ8M5wX+usZ5bF9ONOUl/xH0Zk
+xwSSnoHiHqDS1aT7aR1TBI35s7tov3ZJwBTeQ6ZgTg4qgnj3ARJfz0GuW8DpK7zTSNqfjX5auE5
YtALStkYqfPRMQjez1yREQxymnkipiZ0pX2J6WHEynQbnMN9n7jwTDetLEd6EqNZcGGgY3CIv5ZN
xyvaFrwr1eL/RFiBIYVlsFwKtVwWNjbKi3kpQvUfxZXZB8VFpy1UgritwK2HO4Mk6ykYT3owdeYa
69CjkQZ/6k/Q+V4zU1IOrV+WK9+5tBMXdefFCDJbIMb5xM9tfzOqYxC1u3UHtNz6d+yDOJCDiRXf
3dnDeLmg79Ke3KeIE7VTwR3b3SCSaVQKTL2oLMLYqQA05CJA5FXfNOZPzFJDm9LBWFqs/pE9D2rw
rR8VTy6X06AJf2VQpZqiMAexRqL13hnN7Mein15Ii1qU095sMWEZZhWv528l4u5vmKdNvDYFuGHa
HX5fEQVPRLsi44vaOLgfblAdpI72o2IcbMUZZW1eyE2NTxPvzAzgQlXt4TATwGy29tfqCm9iHKeu
2UQDaK0lZFfGM+qdS83ZLr71k+w34Mr/e/qBjCnZaA+2RhVk+QdOc5CyjfeV02JRfT9CrTG1JDGp
CU5bTYj2J2QDVVA8vcTpBPNBH94UxQEXOtwxC8NCo1pP0iuP7Ix4NVcWd3fWYY8VuIxK3Xe0XjZB
+1Ibo/5g6VFs7a/yRwi0qBvOaaeZuCkWLGojGraEHj5tX/9BTVZAJOPXdQQEt4PEnirstuPsx8r3
3SvFO5QEPtR2m+R1KwGNYpcY7FF6nxn6K97vMb0Y5fZO+p4zPH6AOn90Y/1xUYX7H171ynhDIQz9
qeqhlX0SVyI9p9NXNdB//RG3a8F0dTDQ3d4fQ+ejEOThZjG6lb6MlevjDnYnMDO5AIYuGx44qImj
MXb6xflCZGvhocE3QKaIANsEZt24reqHbgMHpyzT4Qb8T04DzTfgg3NNJYoPx9+cdRoxrkQW/vd1
IFJJQlvjSd1Zb2XkF5jLkaRJlj7sHHGXtGvj64u+VP/C3n+fihw6XaS/RUZvoagJ4e88AEEMA/af
TT2iaECUbpiMR0cF+ZwufD2x4Hu1FVEhDQIQYYiD3u5/7Z8zLQVEDqNB7HnWuoswFqbj2bXn87U6
w3MO1HxYz6vvp9BKFQwbKu0v1Pxw2qygZm2akWW1OrZgCemwMnt2XZ0f+R98rMvQMojD32TqnNkN
GwDd1maB3rlY1fem9Id39VDxobIydgx6lZ8rszfNxjxdJyCK5vQVfHRlIiQ67v8UNfvQdd4eM0GB
Ft2C3Znbw9cD4+HLcMADsbYMsgVq4S0VMJXWJj4D1Vk7JTTCD5MYrbsRejGGwr2IKqOI8d7DlCL+
C6iKk+amzI2aiuz2VlSuBobpA1gvxOh2Wht8B3LOoHRTgpte3ilcM51l0hYNVrmP3tw/22joUWRM
gnqihXU9BAbGgcUWnb0rscvbi/cYsZrIH0oPU6ibBXedF7xhhCplEXNfTrgqkHcVouCAdFWZhqjU
mmfXnrBSmDWZeaZ48RgCnvayjIQYqyHeURpQXJwMm5lk8xMOx+EPLAMnTczhAfplBQRmvs5VlxaC
lRKVdrlEr7B2y3F82v6KDcQaSHgva5R9BCep30QiNR49yiQwgzFTFfYatm/tqrOhak7YJ1T3hXUm
UrK6pzHMDTQCju+8fkD4wQ6pRP9iNpZa5qOpTkEyeRDJiQOVorr3A7kmSov9ymnvVoNvgGRi2Pi1
jC9LvLOFATpQ4dp7pbLk4btUpRlwZRmM2xGy94k/QC+ywsw7LOva3pOSXapBBoy4PnHwbD5JVapV
EzMoA9jtSeoh6mX82IcAs63LY7JhJogQqi7JTJdbYCUVlfgDtxKlxOl+c1iM9474TBOqImU4hOhy
z8FyGVJWucYQnJfPXiOXvIk6IzV6fTK0e7RKLpGNVdQZ7gcXMfg0zvxIwzcVynxpgAZLhGm6UxLZ
bmvCvOEQl8M5+nw3eQpGAi6oirtWWjxkHGYMnrre/7lBpDwVJfiHbUOs8ef6nmvw05Wm8oB1ZBtf
XangulTPO05wtFSKIW6BI2e00NxttFAXCY17e2nJgH5jUaweZsVebHo4qiRE2w2WfnCdOO9my/mS
3+uPJrEoUPlDo1BonRbSao72kda69JORuS+Bo/zckuPZ7H6xbxlut+kuuLn0LpOA9DRdiEY6Mitj
eixNTY7KUtZADK0iJQTs+C0hPOD6ZyCRVucMaa9kTJYzh6Zez7zkXAhmRV05VsCXzeEmVPzusHfx
tBBeQch730E0wexQb45mdbcD2TScMO0TwQJrcjQ9xKOnosUE9wx8COIQRU2b/+j08ri9qL95VOId
kox9BVKLRv5V76cTcTNiHh8CwjAngdk6Rn3Dz9fLWn8gZ69LxXa9dmo0j9+w1lVwbCks2mAtWON4
ZmiW6HyIBlRqhHDZ4trN0wScA/tDgvI8jYomYzJHGz8ihSE7z8ili94bZSpstTr/teK4e39cWx5+
aAAG/4B7B5ykWWjsepQ0b81oNREgxQxSOkBuhRbhw3a3rqlI5TuJNAGsgI5hyhmjM5j/So1b5MDE
nPG5b9U04RmoLTI9OXizQ2QxV3bR4wOn+oGlIGGa6ifW1AA53mchwJnsJt/vdc66Ykn6qMmhwFlu
lv9bHjgiKqjQQHrVCDR19RJnqk0cq9fLsotfBlnIpmPVeCQooF54IQn9/ZLjfKrtE0tmv4zXu8xu
a7tmoK8mPePkK39lOBvjeUmgYxUX+A2BDfJDotw2z6b8PfWphpPrmKuKFDdk8Bx9mWkaT7BX0asd
NXOsnAVFTP+Tss2ILboINs+tIuTfJCWQnzyhYNSZBsn6R3W+4RhltfCi4saxD1RjHIWQ2dkTtc9x
YDP2JOIoICbLCYg0mrf+Xhp4a3pSnwQJbvMbh82c9sTIM5IIukSd2ra5j0Nvr4bedQNQGLQq4iQ6
1yPE+s2aqjM3GfeVu4/FQp1cX6nAQS3LbyQA+WGAP/HzumFDov7W1LVw2STSGSwegzYGGMJqUp7X
OBdF3TplS55nybG++LyZhJrIQBgiWhlG/qMfXIqTUKx54MO/5kyKw0ptEKLZwWEH31ImSxS0pkc5
14wyx6GU4IZzsqrCRklxse0anqK9Gafm/7uecNR2678YspPVtQy2Nkk33HjZNlK3G7hPiaK7SCca
g1A+v9uk83vWRW7nGimaAY9d2QYLSa0cNGzeyRrnPcYGZUaDSHuZ2+nKiZaKJqJ16SDd5EP90PBb
H88dDx78UTTm5+HDIKF0dEuRs863FiMyWk9kgrMlriK/jcGkZGJM25qVJFiOeXwdhCVOW9CnSLxm
CEQps0qEw+7CzHDYlS6zwBR1XGVRME0ymiSV1D7LAzFOK7+KWetVmT+Z1c1gTsYsCCI+kJ0W0y7f
WSPuq2jpWY4NXmqZNlPiBuqy+Q2NQDL9qbuAarx7SBT5tjezGS6WKl9PppTQDgMrua1So2ITXo1r
Wny4z0PQ3suOnATdzbSmqJZRY6MloXatFPhXZj75oewVBPGtQKEQlRqy2yd8F9zAhGtlK05et8IE
HjFfB0bYM9uu3RE9XpVWAigCAjK5mahGU9plW6jmpsibffvpgi+mUKSpmfl/CjDmHV98wK/dFKgq
KE7sabYkN4HPd/YMlxymnjIjzHWbddKQHkRM4v+gln6OoAPImjvRpyVMzHgoan5i5PuWjspG1BpS
r4jzmnsJ+6t2pyPCgYnR7iBfw9fcLjTdZG8Mpn4+aVrq8QcRaPBWmqp9/gjq3I8uCJe5Q+CQOdG+
4kD/ZSIbQg6Oibbib/205ohmcNIY+ctQACEIiVnfcPEyBVMtRtfenBcSjeIsFx89nVcxbXi52D0o
VmgpUuqc4PiFgaqFZxf3ZTFEoazXc3uPowqncek522f1vf8BHEFNHtRXXiNiw96PhsTzjMnzQGue
XeGmlwuDuhMnWT4FB5IuyZu+SJOZejIN/xtBHtM6RuBeFO3aga8HU2O9S9ncXPc7iceuoXNJaI21
HuULsDqK2tIIVEx850ixUsxAhKV/RaI9f2200G/Q+gDzge1FjKZ9az7RZlt2r0IXcigN8J5ltCuM
/oyIgxveLqY9WXNv9snU7GJei7dQen2WssRWODQuboOVje5XYEbRtbUPiEMVZ6Il4le6ugyEcI1d
QpYCNU90Wh7XCQKcDokjagYYeJDGWr/8HJqDhrZiSomNYmNlGEI7YYO0VLRtakDvd5qCX5+t+maX
XOjWBQnR+w45JAwMgC5JO/eQxeakLPLzMKpcK4eGnAlXeULRB7awgp4w+p9atoQKxA07c4I4VAk+
4yMuDA01ZDuvB267NnsxwfmYAlNt9/L5/0RbmsxOuLFGkZSAQf2iykR512jta50q/sHOHeAuHjMS
QDoUtLNH8FlhrXd+kudpvHy6tkNQOB9WZTDVn5jAqJ4sgXh7yvRE5zStGibbOnIedvbripopzN7x
Z2nuJgysHHs+0J8m0a1qs9rN5E+cBBXFpWezZ/UC3rNMmma+zep8GTl66rm8UePxoGDZ7oRUQ+j4
zA5pt/DnvA9Yn8wNjpdvxldn5S/X+Gh9p21SOF6a5AEUEq8/Otj2uucizGbAy5wH/6xuJPMAsKLW
8TiKGWOkHbIL7JhBKDdBQkN9srw889Y3KKf9Brf2eMWANSkzVYU3KY1/TRU853RtLjB3riBhEN2w
fBH/1wKSg7sgzb0jOkz7YA6u/tGd5izg4HJ4VHuzUeWFNNy+SXv0sK2CtjtgqVTxar3sZvPpJBAm
rpNyO9DAVzYEoGQGh/d9fiMHiT0H4hZKIBfrxV13jC8AZgBrZSno5sQfAspR2W5HsC/6QWtwN9dF
wEtps+Va238NqNBIn5cSFGlSoXtRDwKSXsbkqljiZwtfxdjVS1wM86bQ5tF1JQs74QK7EjBpHFV+
XgbIDoalAxCMFedxIou/3cwnW8AawdO1gZqKwS5H4deQmU6XgEwd+3RkSEcHTWd4dATnIMLWWhRY
Ba2EsPeT2f3sPV/muyPruJap2q0zECU7cK0MgdrEH0gTt1YT5AN8p8zo7OyI4CpW7u/O0jr+UEbY
uspRQFhaQp9PkMziW3ZX1mFp6GqTqxoEjLpLXR2+LENWizHWAusc5CBewWcTV0nX5f6r+CKGCN+Q
fRaIHOm2aBeg/8YOjltH/OSmczU3e2NvHY91gPYyWxWGUOoWAiA2qC1QCQz11/E8C8wSKXcVS5Gi
ZgwuCSKFtNkdlbpddtFU37yDxdSCP2btkaR8xmAB/vK/tXAh1ib7jBFsyL2aXkaPhVc/nVxOnpuv
2rX98Wfdgbi1PcBKHZ7vYCYUADzNt26PXdLHq0LGOnniy5Xj4469ndl3enx4qGL9YRc/dCKD2LyK
AhapI6+WQHO6u/IceGEhm+vRI6ZmIBcEvatEkN/5WhcyOFEHYV5KohcLU/b2ZIPKFrp4r7ucvjS1
tT94czPA9V446FsI8vRaoej7zhfA6tJVtVpkPChOW3DQZgTq/DwuCzzE3/F/DXjL09HBthzsSJUC
JpFLMpmyl5KP+SMUDF/1s6dUTdVlT8Y90R12jo6NtQy91pxWcXLrld8U1V3oUpT+6Q1hiMv/yIrK
k3C3pprhppKk7o7G88kZplqfG+TrdrGu8Ujq2iPqY0VQ+CHhQUqgK3aZGaGWu1coozQXEdoqSjmC
roWP1XMAl96mqEpqjveZu9Ybq+kCInxmrmmtlMIW+ejJghIYtFpyHAXehk56qmbLWVwkZqxsJyn+
KcftXWEUBGVlCpqixTFiRq0h04xvZ4ncX5quOO5+ex39mvgHRxN/4o5wH1cAePmlVZrXVD4qB6Cq
gvWtON7Py8N4kN1A65iUrB0xTYDeCWuTY4QHzthAnT7ycK+zYZA8ftfy8BUeAQ/7FOi/kzj/fqst
dpbZmltOCkVFwFQ6veCZREMGmiDAUXGk2xdxKDP1HUDXBZDOEb6KNtkCvBdqos8u1W5rD9ZPYTok
4F9Zm9hx8YW2B8mS26B/Smcv95va9yEb4nksCYQGj2UkNiVb6LiQ3Bp3bneKfuC+kFvfw2/rO3VX
VD0rQ72zcqgCdi5IGMvrYNjYEyzAQEthu8+Pi8y8u7LGvT0IforWZ0IQhtGPDrHUW3wWRyyUbHog
Tn7AqtU8m+oqZoh1h4ZEZmo5fKd8y21LTsQGtsC3s0A36NQnJ2hdS2Q6/jawOltgW3CfkONo7JRf
aeH2RBRHVp9GlIZ2uqhBr7YtqYz21QeoF2ba17k599M8zg/MitipuaCsMWgGeaD7b9vs9E0s9thJ
mXxCxR/8XSSoFR9bc8/1Ufeo5qnGGuyhP99j+vOfQP0mQVg/pJEZl2nkGxvAGjBXx3R3pxz3aoPl
ybVFFlmPDisIBDdtmoaLUwTGB61/3I4syyr8nSxVy11EwVWk0ukmEkZtUb+1QyEvuYP5qXhRA6aM
IwT1cbLJGSN6w0XKpEJZsB4BKh4z2TsjMx7mjnvuzdeLNOWei3Vtwuy1QPlaSJKwQuyi2ak//NZ+
LMqPB/qjVpQ1lxvMZny43uzIwbb3ZJpRQjsugu3unPLF8k6YmBA5fLNJ7u3DRiXfC1aONwW+WqAa
tIA1jyEDsrNYnl9odmeLa+GmWc4DUyxd5iZkPVcvy8OV+7D8rBK7Hzb1EalfesSemcmRo6dW/3Tl
d2SZJJRVsKyiApu6lFNTaWMJfLpO1Rnn0V83XQ5cMubPSsXTCyH/QFWXvMCP2qR70qKqOJN7O734
/MseZcFPJOx83IUP5xTSmjde3YQDsIm8M0UplraHQdaoMnjfnM0GtCHInOMx3RJyiGfqOQbfo1Fl
srN5K5U5+jfblpabPqWdeopGObU5rNsIb/sgMuAlcXl2nKSfgnTCnnM8iPAFAJp4f5conn90PUVy
Q4CUBi3dvcywswJPz0AWcbrds0HHkJ+xnnHZx7LicffHff7TXW8eihfdx59oZ/oomTTfjx/mvsbG
5ZmeviKQLIS28gbqWv6dpeI8f8//M5B+XnajkqXNj8a9JXiCYJH7JtZxHQAIRwdBlGRgRghe/GaL
gnrwRaQIfskuh1sU72BU5bqNhXA7aN0wUv8wmy0aRZOyHy9WiVegk4r+s9Yr8KPF4mDrVwK9WaU9
/ttB3KLCe58wholnZM/vpve6XMn/sL5spr7OPNydB4ekhEWVWSc4N8E129QV4BtREtV+JwPfbKO5
v0JXYGA7K8peUK3OmfMJhVpb6giwheJ/PB1uZvBYGiC9jw7bnR3ybm8uzgLVDNl7ac+OYGajx4iH
GsA+9j96bURVMk6Q/UcCAM1ZjW7e1WTh8KhlUBoUx4BHMa4eoDynHP2fZRlzNhjgTawVwgecRTMD
3N0hiabXZgb4Rsa+D7AHiAdd/s60diQ5hscttVbV2PRjWzt59YEzF4tbLst1XO5vECen71/pMi6U
5G8VqzC4ZhcLEAfwmqyrqaR+R+hkoEO2ITuUw4lOkpLThva55D/c16fthb7am9kJCfwJA/oBoEZW
aumLoRHvnL8HKaQbI9f+MFzetRsRd5NGZjSvbCw4vqadYVaguXeg1DLuClmE/INxnKvb1QVzJzSs
iGGjBV9cD4jK+b0udLIcrXz/Wi0eUkjgvrM2zwbrwnOiafUe6PydcUzgRS9fMxx/JrhOZnteh2AK
ztvGiIqfDBquSbPHs+UYIqt0sq0Cjqf+zRw49HBCvPLbh2EI2jAKjMCKtl7eNgmGcTbhWtSIr7zs
fSj2AzLAAhJPO9p74mEW7A9GxM+ir04IqrWQf4v0Om6hBTj3Wbcna/MitiBiOkuNMXQ9NwM7nH4z
WUKELHdrivGQhQCA0YYvmBnEux2LS2HxQHBdWU6YUkHU7swQp/3a0roj+W0HqG4F363piG/SFgfE
3uFWDgzmDaWC4ko1/fK52POaACfB+0zdGlxTsOv/VKLjyFUSaHHTzL6f/PPPH7iOkewUto1kV3Fx
h4ej+MA4bpPkv/qAFV2cK/fwQ9BOUU+iyoxYJIdSONRp0qFSWProDvNViY4cQrXS7oFzqWl56gd+
1rxk8TbQMaiC0nY8hdL2ebeiUdWN60TZiRkx7M/ZKNHSCzZH6Sf4o0YDc+YvB2OnWV1ZqeTAsHrF
s30tWaMuipc0BjUsRdN6XBMRpYag4wkbwUmeKxh6xEAy/1iQsLhLtE7el7DQoyEqsn/9J7J8adcC
iu8yoET0QvIbdfBuaYQrasgBXNi5jqaV4IXO3UuuxsNAakw9XeCjNtrXKNByYttJ4nNFR/vD8Mwd
eFBYmagVGazn6+xSBGi2Yebtk86ywuOLkpgFfkyipDwADE9240o19hoA/I4FEim6e0sYa5zbFVio
UJfugIPfjc0sMsww4wAnaTwrVZqReuzBNHuTtIdmknOZD5BP8OZsYagOKmO8xGFpb7I6rZXLupse
zoDnvDmzSuzdtiDUD1axKDrGNkjR1jNvbu9ZGHE0gwpxhhF7khTrSuQFTPZ6r4c6q41alqoPWLp1
4IEqWSih0Sy/iA68hJKbx/HlpuSzFK8TG2cJm/GTJd9KseGXpuAS14CyGKA9PUajTNukw+bPqwqz
nIKXIy/FHwAO6/HJngZq0cKGnGEHdGixuqJofKSR1XPTaePqeyVseBbZVrLofdXU8QdGA0X02Gr6
dFHeuMpm44iCznHCtn1sBR17euI4L/3ZNVPMgCbUITLl+63PAq0y5dFZSllyxSx3KEMbCiHNcACM
NKkKYRxcTIv4DCC0YGD4oopY8XIIJG4+xG6tlEgf0WPWKGrvAog67T3U7B2f5lcdOTc8A5Ip1/Mt
pOW4NpRakOBuc0PbdA51l1xL3DRS7cDTYeUfKc/zKHLwwl0eap7GdNlTKQwoxYnhg9uq7lY2D2Ds
QD/GAlfkO6PgIumDmT2aqw2W01AUZbV+LA0MlfPYZH+/yQ7eD/FeGY6jrvA8ZRJ/7cxDEI1kmMum
tgLUAOm6d9UROe8Agr+DyORqSgVLBjMvGkCfo5EPWo3a7syRwhy4Zq2pNG/nWjFnwjYXrNGjcq6j
lplfPncOCCiRzQnd/wDmoYWu8JXZICi9tItiN5AJFfvEbXJy6c3stOLGcmjJYvlLYY7KBc0wI8Uw
a+AouV9GpE2SzoS1M9IvFHd9MD6WLLYzX3TOwDSOVi0Ff9lqctZBgLevDsbruSg3hoTmx7lnSC0g
cEeOTRfxoUnzY+FnOYfWHJiZDmMajIUnKY+naTBGyxIvDZX5XDbXkrIG5YePv/stpq0EZXK7A1I9
L2DPLLXnozHGUYSnDF5s2iTx9rCZNztHy5p64TClIkeQCRBVmxEsLM5J13Pb/Ddp7pEVOg4KU31l
V+dDwE3kiwdq7XxjzQZgLzo6qDiBODgF5u0ba3Kif9hCgB9BOaZYjsa22ZrAMIn/vw5DKep36byT
f1FyGVOB/HBClCsihIA6lCh5t7ovjIRnQHiQmbBJ4y4T2RVmtKzrDDInPdFT6goRvKdYwSNkV0Fs
xlXk7LTMV0ituCt/4U3p8YkMqfXxxCHDlABTCyHiT5OBSvEWNVZ7rx7z/YNfoCRwOr1OcOrLmoy/
V6V0567wK/b9wA/QIijCdJcMPlygEsRb9j0IJ7q3MvDFKshsy2H9mwH41GgFAOgy4dTYnZDvDHUw
U35dHtcmzW18rKfOUZC7uC1CxYNX7AhVblgoF2Sok0VlY2UZ3L9Wu+yTs2oLcPPY5+4Zh3wqvWLV
UG9H0whrUX+wp2f039W8Zf16xjXqJHJQ2grWU+8I0ux0FQhujq+gA1JpcHsHTIRcy8GBw7c5DC2f
jb6aUfKOjF1SiE4WhHBZ5fS2TIZH3Q5BEPer4Jp8y9FfIjeE8wSFMcpz+7VOP6Ua9RP+VggEMI48
Zplmb3EFGwx2/Uhjf045Q4MPr/mi0OblUgv68HEbSS4L0BWy3EXjGYtTMb1/ob2LjzdoN9PSeGm0
bxnnlkr5g6ilBV7oNCt6uVSQpR7vCpv7ZdTLUkRoqaKHWSBkQ5O/ca5JDjsfhkPWIFqCsxN2++TC
GXFotYnI3RpbFvZInuY+Cdms1ne2TawPN+xXwJ6MRzxFr+djKJbvMzwiuTD42gv3JcgMDt9Gojfs
+9V8UlEaVySTPZPSlQxn9FLmV/hxlqaJXFQWkps2GSx6kFSBy505aW1K0tIoa8j/NI0F8pbhKw2B
JzpABgj3o+fk02DbB1QZ7xPLzbzVuDCaMk9O1RKysbSx/nlEZHjWyNK7vCI464FvnySas165SZXu
/ocFePgH6xRDducdpfLd/VsD4ntTxwT/X08GL3rWZZyPyeA+sBkTP4sDzeKbLP9hnvmb6+UOEzgr
mdiUd01caZWRPHL2yFl18oBD6jE7omlAHi+srpKMPVhqVbL2iS0L8erYIYnmYDgEOrntnV5JToVD
+c5RUmDbBcu4CO7nHYMYfxZqiKOpdO0ZwhAGqu+FOxAKJUUCm04K3GYYZa3cZanL2emq33hOSAwI
Kn43hPHlAAAc/QDpynGQHHhunhIGYbmdKZ+D0vnw5ygq5n/u0IlfDLZM5HA2W3bbcxeC6PkmoHyi
1xNrHBW5bGFlKDJh6wFnEELH/7s+zL4sH0cUJKbaLqRRhDlHbVRCwcvl8w7Qa5wQdQyc7umDWfQl
mzQolsRBSRHRzFyURghASZ3yK+XhI/bIyl5pGk/6QAB4gNObtQg4+ZXPHu47YXDrlp4I1tn+mb7d
+Jr5dfCt7hdOommaBdb0TC5crfKaftZtfG962t44yBAYHt68p36xi7nQN/LivBFsiVjWDdFMsB94
TDgAkVrech+lrl4hfTx/rwNRpnVzPs8vp6I5ESP0Z/DqbXp32Z/5qpvq9Fr47LkBzMFBsnZpVb3u
KvdstJmkQaqgNEgRJc6i1Y/Uc0qJb7adP/JkyS/cMjS60cFFHWYMywDXLNFiBfeSFbdWClerZyXJ
D/CFHrKY/9G2mQcfFjQlrcjT+QciP5oIZu2Pfo53NABQse4yzqvFEWa4EYJhf0YJaeacsS//gfMd
yjlIWjJZ6pXM/E1FaZ3Az6O9pXc6iKzNix5OdtUPrBLRTwLJkoj3YpCfV7vBvziGZvz2uS41izQ+
zIUd/xOIOlEdBC9X6Gn1nppoYHJW4/AWGkaMdNGSw0nhTbdPYT4TZ6rGpX82IuOZ/1U+ddE/aqTe
gLtDSBAJyWJj93NoW2/kzkHq8WPFpdPqKO4sOvlJuKVZDMfuVGWwpkagEOdlY3ZrfW4suInJ7p3k
d1XeI+2kspqC+p8IyGm8JXlkMfZX4EQN35AdvfXqtH9DMxPTRkMq2rZ9XCl4RXnicbFQQLrBCelr
6mZ1amDVRVmysLWam5vyuDfewnYatDfOyGrh9RSXPBd7akMAPfu8LoFZ+VPB36eM2RaYSd3TxkXQ
d0ItZUKxZdiA1e4otBc+3iMd0eqiR30DXoyL38YS9PrpsTQhlLnywj5hdQm4dwlZk1khQfBND/aP
RtoXKbQeg6qfjipGYuyAxFw9GYIUbB8p5wDPRtTJxDZHdrVe4aUkNBece0/QlUh/MOVMJQb0BoOy
jntZzAcMcI0Y2Jdra/IU+fswgtfVZw70gxXgpeRyWTSLZx7fPF29uw9EhgmgOhy70TP75z3AHg0l
21wTzf/7VDdxJ+nGvunxdK/qtRSN4BHycmNW4/NIT81Kshzn9vAA3ecc4Fc0stg++1y/amQbB+6/
pYO8YwxPWzVAFcZJ8zYwXJoGQ652g9h9GkbCCToTVGdpsGNp8/mI10sxpATp5w7GzoyTp5IpilXI
c7rSibKDJwKewGR5TdLkbd4xy7dHqSQ83ImxRMXxwtPZa5tX+1cge5mSsGtdu5h0eT5Q5nGu9UIL
KbAaODqn+yd/+W6qWid1K6jgjgJlaXIqbmIsBUrKxqw/MT0dUo4mlt6qDYofiMnYbrJ+Pt+4zJHM
YhC+NIFEt6xRtYjsik6p2iXc1E0V7kSWm2rflTpFh1zPoxe5xuiDeO4+d3WdcqeME1ISPq8HjcpI
BIbK61nNVK32wS5QNLGbqX1pVwj84ZV6iXtt3KlfQ9fu2jj7Injdiow8u1hKGBA34R1i0VkYhTyt
NXHOQKfRLau42abNVQcXGHVqK6xyUI7TiTON4eDDKZ0yhCcY/wn8dDHihF0w7f4j1MB3SbdDizAR
f96vDW8BaFbNAD4w0qwxrzcv6+sCQZSzcDssXhR1FjHv9jE0vsVZ1tJomyn1BpVK9OmDskur2JAj
NqdF0wtjvpl64TG32s9+e+5nMCqyWJy7seH8zUQYhAVoRkSRVNcS0tkirBfIboKgG4g6eyVlqDRW
a5SJA175YK/GWOJ5WQGeq+6+2omIpZ/mbKGIev9zZ0BKuyZdDV7z7gSrwqTi0ZRYqA3uvTFBadrd
rWaW4EAD37UXIHASxnDTTdh0FgPNJzE+hoeLq6L2M4UcU1V/MVApnMNczooE/u5iAtFxZfZmnDyC
KAnDPhuwRlT3FsO+Xg3s+r2UvcDNkVO1WIGYmL9+wHyeCumXm9DIJWRQykjSbjVwZHJ2KqIDQ1uL
qvrxFbEepW2wqQovVVrymKmkUreNE+L/styWvEc8/0wyu9SsOUZFWjkPuQV2teCviTxam7ABIY+n
s6YPXkQvNuqZz6omNMEwUMuzAVohtCtWFqfsRHU5v09+V5KXIAIi7MvaaC7CTSh963ywvj/oX7QW
6PZ3+j23aFErFI1bZgeKWWaYkLgcxeF67MwJfz+Oj0aLwDLVd+tzCN99GVD2nRZlPzmtTHWyqWAJ
ouJhHySPm4BEnFlelCn4c3ewrs2eZSVk+9r7DjPrWBJdSkcYrb4S8bE25Bsw01/zuEzknpNIbY00
YfuoSDpuCAZNGik6BVPj+/0YSnUCMNfPGntyxGeU+MOOg4vw2t4unXQFg6h6/MLwen/W0LZ1rIT0
tb2b+tYqWRjLl3Eg7jpVZUmUerbWrqE65XY7QscTcya8qDaW8tPzTUeNoPvF1N9pdeP1WmDDKfau
qGhZS6OXZiJE9/5tu/8+CcWI5SvJMXF2ElUKf2Wvr5jq/H4mrqLKN0UHU1dcAoo6JnTaMHpOkGCD
bVNrhZE78GjII3RIwrsvguWUb/qlJOvkrqwfaw10DUDLtLO6Y5sCZxdywKFmAkRoO37R5HR2xXh0
DRKIPy6NvfoEe7eZcAU0gwzx4SB8XNnFB6msrlcyREBmHmK+AbAl+OS+NuR2MrnUMFGe0oT5McDS
zcKq1H4yTCIlpHsKBrIDWHgb0UBXAHt/gi2PB/89O/7uff+cI7ZsY9OYpgOVVrpFJBwu2+TdoCb+
Kze7nwOBWQiLCEMwsu7EzDeCQ0OaaI8pNQZerKKMNMDVBlKlTdacg3jiNx6FSarObCj6G8YdHUqR
boheR+5fgT5bHYlbIR9WnwVm9IlrkmoOIdHXPVRtAN93XNRiPvKM0EC0BJ31cNwhVLbyNBUBzKLB
ig99AVYcZXwxWYOUHALswU1JUZfjjpUJpOpG/JHe9Hy0wN3PHg+i6sjVsYXLrkgNNLix5u4yzJP9
CuPcrxj8Phmxk4FndXHrB2pZTUqZd15J1fYIotOLFXavZlNhNvlGCpAYe1vBRsLcT0GaiMwuEaZw
+UKrSPBugg2AunxJSp3Dpz6IKoVjYV6n86qn9nVbEPMADc54rcj5cy8U3j/2yE4yH98VICEgHvC3
Xg0yUprmwUARFRcs8rtrht3EEiCPI3iHIvXBvxWzyH3FsDce9thARhL43EKyn+uRpBt1pvLL6TJi
tfBILWbq5saOO8qUI8PaX2aHzjxak9OGPB3JFFPQgwxN2n0dxnyN80mIvHM+3oUb/tZ4UAPWA445
6q3AKQxLfHcbotJ+AabCj8FV/dGJeVey+qj2A5dCA98MqOcF5KoGxFeMW00/Ss5Ja0H8A3jLyqFb
Py8/issHWpOGYp4iwiBLtH5i65xBO3iHfXgGbirBPoa5eWn7scrY05CRMFuf/37WCoJtO9xSYLTS
SLYqhmQeTpa+Ltut1KUj0DFISdxjeH5Sz6wMum25PkmaPPz2rfPsU07bQFtjhUL5aV+YhqCQ/aNo
OR62eyaxGCM9jTaJT1Vc+3sW0ubD4gfabgynrC2G7n7Gc//odxGFH1MTilcd4hclNUrQPaDNwtEg
UGlDnDMIjHbrjLB+aEnJtWdbLwH3R7laq+YzmkJV2lWGwjNOyvdCZ5G8hwPyVewl+sxVz2ziO0xr
fWmUzAfEFc4w/yNg4GDwPedMx/sDQCk/1c50nLGtrbL8IMlyoJgO+j+l74mK3tA5YXitazh4Dmrb
PnZYUBt1mTCY8tXKYx/efkePrnE5GueUP5S+0GXh+1PStmtmOR+rZ+X3Z0AswV07WghsE9Nl2k+D
M1gfwzPxiDZBOUDgrmExjopdPotizaSStUnwZGY7n+Dirm/k9HOPb25HS/fsbGa6gqmJA/EALRtA
APV1F2TzdrorxK/0+iPIw/lJNvjFnti/3SK6XBoS2va/jqgQY+2+0RFmLRd0v77u8X8ANIuLG9FC
18Gjvy11BCvugySBV0Na1PjNf25deU2HeRDzSgwdmtuKc3Y1rgCM3/AC9oVLBhPzWCkTu8OrKpWJ
LhqMFdlKVU09SyOP3ikSBFuaRtCaDzRQcjsFZppFK0o3TjlpvZTJ7OXfPbwXK7VRXcFwpphXFnSh
NvEZW++Vke6JxQfRivG27lw+FMLsP5lk2x0AZXvZwN5LdakQz6+hMqnym2a5eykCjzFtSYvueH1s
TioYzH21918/MZPo50oHccb7G3Tdvq5q95zi5A2D+AbMo96GRv5b4JTK/hCz5e190VT9MPgQ3iNf
sY2LEeWCYHASRkQ6TMC7y989xMo00QwDZxT/yOO83Q2NfG/vKgadLbIloz4hfD95/9DeMoG8HyfX
UhRt4eJyBgqE8EwCOq+a1UFLqf1dvstnSBBm5+ae4NLAx0F5OtbpMJyppRhmVnLkpWFHXCGjnfUI
MC9rUo65jCZLJouclUAhFHNQQiU5GTKIL11XZBPfnZJoZCIXhGHP+088866jV2vhOZbyKZL6wihY
EK83TNkIA+ZeS+vbCQQ7fWNtmzNiqZ/VsrrsGkxKvjx2wBmbzsA19UGKSDRGwAPWxboHVHQL9Phc
BzO1y/zn1jS9eZXhcLrMvPBlYXa+DECMvuh1x43wUDjR2q5wDVG+YOSb5OuIDuPH7fahUdl5WoTD
Eu1sliBZa1+amdcYUKkI5E6X8lqFuYhtF2T6Js/KkIa5iZ6MYq2ZQB8D1268XSZ23GG9BkJnzCqg
uRlo5Z1btbmXicHvrw57SbI4xX4roqUoO9SR/976cI8z5AotFTXrAG+wAzyx2piroOIBST+wTdLy
AYtU2sOiGkxpI+pRcEIDa3Tx9XDRUEDp+Iexm2EwAdvZ2IyMRNV/hefhL6bSrgXFT0Wt4uVOO07j
p8zRKSmukrfXfjLDLK0nMdzFM58a/bnDdqeZ7GmEy8eFMgUJnY91laQywbOzJru2RRtxhj1u2dFz
63EGqG4nSczV1Hssv14QajdYDVddCtcu4GYZcl74Fa81E+QaTfRmntwdc6ll6ISHbiOhz8hgpM4H
tERNJxGXsVizE0W+qMajt7bhWtWdDbzSGKi+LSWbxUKaM5v2tdf2BvYalq2QP7fXennJ+WjCWjIc
ujdAmKP5f8JJlC0X7Y+W1AJs5UOe0jRSTRflE1A6uDowUI9CYk0MqZlM01WnSl0VKjnJpdmX79Cd
V+igKg3TuAR+r6evj/VaDxy1J9PKomq/h0BZLd7ka/PjcNbU6l/ef9FcZTxn4zQP+I3SfFcJwsZ+
OV+fy/Q9yOQKm10G2y/vbq751OaXyRHJ1XGQqrXmdx8QuWy+horANeaQolh/mqYHI1m/Chpq1it/
8ffFomMdfhcoG5b7C33ourBx6f+CU37if1C3KMWT4qoXw018jJuhY23VqM/NsogJLNUpz5jvTnWG
pIS8VWhZFcp6+NY2ysApOa88nEMpK/An8/8qHfjt0gVn+iTThZClLDXmUhsWBCSA45LLQNFRZHJr
+mejUhaMDZnxgfxngZpDGklRANlUOZKfpxiPXtt5iE/hJ3LcUVniCj88MFi4E51ALy9acA5sk54R
ybyGJsGCnM5MD84/bCMWxHlZ0qU+4TiskDYqDZT8ml/0AWO/Gb5NdRFaMVJUX3hKpexB+CUQF+nn
QuuRMN1AvuRmNczXoaK4zaL6uGynQDNB8xNIaAt8ee2k2SPuw2RM24NMN54nkj5mWRVSc//0ngh5
7NA620DoVdFX9xWsiJndSLWX+1Ipo3w6vSgq+Zj/BrZq+xw11ttd6od6edZeuIcoejrqPvXshMhx
42FJGrcoDaEuv8WoaF4a6QksR4Y6/4N6aMYbrMUPcgrkOT7CgF8FBR/CSZN4lLHl9XlCe5ngNXKy
RI2tXO2wLnlZvsBrrpQk1BhicOmC6sG8Rpqfs3gvEAa1KkMdbw2Ar2izqZnKMqM158m+lGaxLxpv
nUGyQ8UvBbPpnqMSTej7CK7GRq++fAc86FGeKwQbHgpZBD2q55Gr52qsRFpPGudb3lSGwaXBGQ5n
yVmg03Bb/TQRHVlndqUSDpUkuXnUGczKLWKXsQ4wD19PUQYnSlgdH7Asn9IVbgr2jjPF+CbxzUkZ
3AtmqYORrKhkBh3GHG4I+X2vWxIkQnMNUBMMrlrVTPVW645N7LzDomwdi9IIPXdkJJ5s/CzePwYT
XejhXBek20aYWK8yzhh4KoY1rMjGioWYklhyVFAOGC1Kqs8R8s950bCOh+II90iEJy98Y1m0PV1Q
rkWiZXbNHHgpQ5kIfJWrC248Ar8U5qpfmuTkND4jSmkERJdR4eR5nfaoquHTfOxuA1fPpZk7b8GH
MwXONzBQUePOs1P1JNRQRPPHwzBmvUSo5ACHNET46LFBRgpJwjJymAenkUkH6pi07Ezzh7X2qs0F
Aiy8uAwewEe98U78k01JEkrJo3vprqzj3nUhCvSwNoQAM8GtCpX2uP3oh3uzvxGHvoexY9eN3Ubp
PEJSvaxsdue/V6N5P8RwiXLHX3iyVeksbATtvnhNQYItW245smpLLcYQijkRw+5jUP3/O+UDRqid
MXlVxGwUDrA+AnmUNwC+sJ0g89W03gDtRWZM+mKqBS1d05YaGnmjh8vCaGle8J2qT1QaAlBt+9D+
vYGxHvbTniNUF45hjyTDCduET+mBviEHuOeaNpRFv4BZB9iGVfo95N4eSVBTfp+2v4hdyUiNGyzH
pK3tZmH19TBMjtQ6fEoInJthyMfxuDyOpx6xxArCPkL8SXxbFfutWsNC2lp9MEZAmsI6XtaSU8zI
03+VU5DsFHaWLTOMu8cYc0DFIp5ro8leKAm+ZcJGV79cQhJWpTo9mGC9YR19cK16MjvqoHxCSqe+
fZEZFDPvNC0me3R4gQ+XHU9/JblSJHSmTKuPehwBmeoorTj9JnIRwQ/JIIW/lZjA2oWoIWkn/eo3
l7rR2o9dW6mSoM6dQM3pguKlSIvkdruv9iUgB57V68xtT5T4P9UxcpxSs7qN1Ov5VV7JSv1rbRnk
BHRUojRYrgn3ccJ15GfxOP8ajNfxwgDqPLp/ySf+d8GavukArlobLTW3w2WG2+D0NASUFdHXg0dp
yW4WD9XRNMMaTi/axOXuPvYVZOHKFRegrLCvyVGL4KLAs1Xh9K8cQi1QuM960fIBUJf6Ygq2ME61
oTg1XQntBE+1EKuMJeUanoEvaTksH2FXC/UvVl3/N+B2d2tUkL2v78XDRBRPXgcxU4K0QZgHBaQm
GbQqz5LIXaltgD25xWShcH5y7Uy9tRYOTswqV6UaOG03ACKTjkdmm9pmTckMtSBCVimsmpARTiTx
9RXtzWGaWnV3cHFkKUOALEbfgyYf9S95aHcPjbaFjvDdPCZOIkUyPhtegGcFykMGOG65+GOkdl6t
xUMqZ0YTo4eRb2rxJX37/HQQgJcizrhRomDKleYBy9TXQIZKjDiSpjyhOGZKEfZnLCv3iihStk4I
1wzuWD3yqcb5T/wpvbrxagtUW39845kLUeEpT4L5lr6EZMGzhA+6m8MRiX7jz+RtinPd+ZeajCdF
RavYeLlBcvHR9u48Dxr8uakbcxO+CtcVtLBqtWB/J7OAkQcjUR2XndF7NqEW45FhzsnfWJ2qvc5d
yskQBdGl5/SnWR8/7kAwKQKaE46pgZtwblstnUk89yJ0H05Z8Q4ewAioJdRKGXD3UWyAVNxO1C08
ibaQJ55caiI186rXcKHPF1ZCtm4RLhITGpFvnwpmMg/39Un6EkZ+GzZP+ymn67COcaPfuKtxnJO7
vqqqgWlTYnS/Z2jx3Lyvq7qeZGLVMwtO1J2Ppp3jLb9i/V0az585WFiLvToN5AgOZN7hFShwe0ar
bmoKDQTQUzqeVjDhc4NmZiFDu5RlgQFkT4Jz57jAq6q51IcsgvEwI5tUYj+cn0+o78CsDSaZtrVD
A1M530Asm/gyVJFO1izI0jqTvMVz0EQLfD/Dr6p0yF4dwWHs2RKQgVRBVcg+zV9hnqajCg6CkBX3
MtBb8uW4M9WGSkyvYUlGvIijWUFl9Kcde/7pc35oVmydbZv0V4bQZ5eku494JHdi1hoopeL0G5j2
zD8PUkCHRASomsEnRnDYx3LEW4DskF6PArqX+ID+dJW9zGyEobMN85UwuJ67pPClIwNv7QMd7aU+
YxGZtA2UsG08CqgO6Vb5fwjO227eL1n9zU7HDTSGnFPuOQS8ki98xdjrvUNEbADR4n0aeeMTtyz8
ONkPX1QpHWFpZnqoEexeNLKTKcVbUE6YMUZjthACruL1+j38TDggkxxUVBjyAxNJmlqTy1c2rmuh
ubefKIRhZWqUadUghBccsEu3gA/kDrwao4weOIVJnQWCJVAGVq+sA62Dfti8g2GJwysiQ4Zqv5Ne
0s5WZuPk69VepZd1nLR+pp10SZpEFtiy5BpMp5PAQ7eta0wJU7j2B6xEvR7Tt9MWHauNc7HF3LvX
8tSlIZ29us/uzlwjWdv9RDlFoMbpYjXeML8Mw8Fr3bKNyp0jHGFC1qJmZ+rO60jFZiMzURYVbmBN
LHYeVnHTu/9sDCRfY/PkYeM+v0YKngxW9YeNDbOiH9qIvCOeBsA6hNN/TSs74h5h18yMm8uhDHqs
Wi1E25v7HndKyodPGXVZ7RRL3RUiWSGipHtDD9fqEUczeE9nfL5E6LrPS3VB4w9WjCDfRxQl5yVN
wo78DSk6KlBH3rakA68QCiyET3AMKBF5UxaJChtcmtK1f1hU1IRHzd3Ql29zG4nJ//aALTe5Qdps
4iKvpVWg8AI+tmkm+rmpsNxsvQmIylcnwxlMeHufqRx0iCYzjqjyBWAIS6/nxGakUo5VEKLYdV4V
EY/4rGuzdFVtpXmcmS3Lahp2dEbX2Bw5J3uzV2Z9yvFdfOPX7QYTJRTZSamtdLPNkcwtQHH7KCjZ
TseKi2cEyFozyjffo+/Hzefz7G1OOlHzWT4mqxkOSOdGRYAXc9TG731HrQg4IMVgaduvF33p5euJ
qjWO+ZoN3EGUP1XEsECUBA/Q6CE1rAPGBqo5HT88dmWLsmdJJXxOQocBTCgVDT8CSKSHvI13KB/F
iqLHKOHnDROuEKnX1UFYCUkfDlQnC8KbFfcMs17RbsNIkxzWCFMnY50T3T5Y7sNQlNVCB12Kde82
OBsN7/V3xzjq/WFJTEXQpOb+Su4CJ78nMVAunhYXoPRPA3pi3i/3A/v9fRKXs/WsTbeU0UB1mE9W
ZSK5jbWv+2WL/Ui6W3Hl8iYwvLveSvxi4dp8uMs1WibVgu8kDmxNjROrgyiZvXCZdUlICaVy0xhV
frobNRIXuAmk03j4zF6TL2Is4QbSQKBC5azTptdL2PtV+72unPuD843pf561S1eJ4yKd8ZOK2/+e
ngk1M3DE4ExtuJo5A9YNAZCw0nBmPasncQogImwSnCc/WZv+5tK6bO1fqA4fsI0SEAEFLHyuwk5o
Xwqpqu7ROB/oDcceF45Qowj4CHp4Ff9IF5sAod2UTbAEcF1CMDT+/jk1nXQJk8CX8GH5sdW1oIhW
YU+ymrlBCy9mVK7M4ECZP3H5QLHnWogLGOfR9pUPbYgqMfbA9v9XzJfsAo1wZQqk8t0WRhWLtVt+
5wpHN+DXGPAMcFyad6gE4pgjvUdY1JfFfZ2S02JxaJgsNkbAsmc7TsdvgC/3L0njMf/8ZcqdcYHR
NnF3SN7u2xxyzRKZBauYQB5vdsv1VuWP65Gjq4L4RI1FYNB91BF6JhElMEEec+Mm6IW2aa86jsfZ
EdSxKcJd+rZuBTGBWNBmC5U8x1Khn2tkstENykw2+PfbMeSmZ8U10V+yO/baNrP7xhJP2uAnNI/L
rKQQuwwKSV1jKALetDFgVxcapIKlhlWcgf93kTfgGdqd36IxhugkmwRYtmqcBrpKkrabnkIII/Kf
Usr4/NhBP3JWV1ro14mDGsfvA0v2w8ODQdiv7msHwXKJSsQmb8TSFotFpLoM9BBiEPWxsW7TRPKm
d8UBVRKegEoDeX/9L4rZkVjnJa052ehNuprfvKlOmPqVZCxD6ex3diW4/SS5OpUeR8ZVmEtdNmFB
6s0I4fYEB1Ems49gspcOWS/6XEOva6tBBRaDc1+itdaqgSMf3HpZ30H9ZjvCzAyybDdYPWjYimsN
fHDUKnSnNHoebAcLRROiZI9V1Y9SNP7XbMp/OQQoAe0Vucpzb1LqcRXQLn1oyzC0yfsHYO8LJn9B
/rWnEXnUfU6iuPi3ml3Tm6OgWgbpA/3umBMvikIi/RI7CQJ//z2NhCb6mTWonTD3/4KBX6nhM/80
GVQDkIyf2p88t/SaJiNwGQYH5jXC3YEqvvfDF1XUtG4K2q6+JDBSHowvPO6Z63txWeDloEgJ6gVx
89wPwA2Hl5tTXjv/cBT5HjGzy2m//8jE+L4V4tai9us6tQWXPFsrBaJVJYpiqQgv3ubBFJmX7hHB
VQBTAPl4q49XB4rltJM7lOVqEZLdNqoEvtCpIQv3J2DYrw31DMOTMzW2WBuZ6Utz0gHt9i4W3xV7
+Sm1a63JojIyEhbek5nblqtWUABbmqAK1q1nYCA6ovpR5wWMKEy+iQx1xQQ18vlkSfBmZdx2Zyj5
iwJylpgQGBMrsH2/dOgflqIrcEWJCYkteHWxWcoE09ADQkaOoqT7hbYr8YjIeVwMjAiYn7adsJSl
DOGWdetZBkzUm1pu5RZyWPu3e9UgWyzn7XfDLFt+8rfqOqG26Z34i/0pel0YhH+t0vCn1k+thNiw
taLXuAnokWw/tR7TQum+SlvrJeLK/uyXD4lvTsuL2MsIA0yJqCsQRdPzLorLm+0cdE7SEcILQp3q
9Rm+POYOXfmbEz/mzWpKMdt7X5BirhIigCkhs21Y8YIVQbgBR22sSkszXSOgxAYn1n2ffMSDoIyC
Tfvfv0JbO/sCW8pEcaT+N3osFf37KsFNsl4RBzmM0c9OdIR6pcbuXA9Fafzyke1ssyH1qLbWy2g6
nr0qg22lLtMumwEThlD3V1/ezlUq7wxzPfVJG7f6Xcu53kgUcJ44z2a6CXINnfYlSJdOCDbFsEWw
CGk+yD1djQQWMCz9HRxSbGULbfU+ZmzcP2yhcjd+cs0tP1+yxnxKAA9ZnnbgFIC0OINOwE83lktE
f2G+Imlk39E+ApCdtKy41TnRbutYOPFMmZvj0CYnQydcQMbvwRtxgPrnm7eYi00BdrA7OovgMsUJ
iRA2lStQ/xHIW2wfUulLtPgw5ZtFprUOkMeE0eLXasCCkIl5JxvHfiY62Bk4HkZA7odPTPf63iiK
jic4DVoIl9V2ldweJ4qn2JWvSyVlAIVaIxcDSUx0DgY3XqDhdT2OjjCflNOerWWjfj+ewJaLyMJH
3cQmGFxgMjtdpwUUnNTOXYXPqj2spkfYpuzKWuvgy2elgcWO/KHH6Ju6SUpfrgP4/To9C6yQjUM5
P/W96/15BqeCBtCtFJKwgInAYvGKNrEDyW6FMRv+GLJcp/574TmSq08DHMpY3EB/d0xIw9hABi21
X8w9beZZdktbMAjz0A0dFBx2Rjs0d+Z0H0h35tbEYGbS6kIRC8RfIcFvaMkonO9BuhDDaSFF4KFi
mPDSLmRCK1o1DkL6mUFyZ89+pV42A6eaeCLRHVAqL6K+VgP4XPFqs7bWyJtYkxhmLiQTUrvytQ7C
Vd0NtwMfWKx7d1HwTRnNMi5SwZBBmlbTMXra9VyHqkIe0EyRgRtJrw836uwkLnbfP/LYvZ4X1Jp2
0LrwiJH80u3LojWCjRbnbUMDyz8px4J0yR/PuGnVvTL1778cUrbW0e7u+7mIrMVF18Lbgr1lrLJk
0OuGMsxk38JU74X0BoaHzCyM+Mm4OKPvEP2eRifVN5J3gC7kAzF2Hwm7d9tQkGC6MTaIBgZuVN2+
zxIBjErsQxZmB3tP0E6bzIn6Ovz5hBSQEkrsYU9IKc3GgxF7ocdMItttJUJ6SL8dOSwr7+4k36SG
83/57HRCnFxu3/g/MP2qSsv2R55ZDCAmmwlCRa6XSrXUycwTh/4yw6u1Rw8AqLcbx9C4jAsljY2t
i/ib2xEBJLPe63HH/v4BJI+fwLwJteGPzwxA4iXzQE3IcdS3OCynfwSBkA1TwSCJpVOLDBKgNCPc
O7MMWKu4cj3O0dG2VIQNMzhhIcqpQRZgixWr6uMuOIG8P5K11/XShjpa54QFaDZNnf51xAwxxF8C
9uL5XE3Un8FCrdfHqx30zGruit40L8DAB4GfZoy1bydgUzaoMwXw8sC9tDpUjEb7EiOjGFA4zbiW
gC1Vsn1288foQ2kU2+Yjwhx/sAApFjItrdZIC2wJ5XetdYKqHyE/CjZ99E1b2ltVezaU6eBr0GDe
YBdGURsoNWfcHqV0J7/5lzRlHMm/5SRmWZro0GpodExEPVaK8z/XxnQN4YwZJODyAZ1LU9W1Ebn9
DQyEg2RnkSCo45yukWEW09dHw+wia0npQk5O484fRBBhRe4scvEdX1CMy5uks85no3BvTC44vfdZ
ImtsqjDiMCb/dfc/g9VasXjU5DA1UhBpOHJ6S/7yGrjq3MaE0cSF4mBMr4X9Sw6QuMla7VfNImx2
GO7S+suP14vG4P82SGtsTySN2hiOnPh4ktxXp3UnUV22m62AREYCtKS0nHYgtcbeNPMVieh86z2w
KB1v2MpqBLHPrP5vdaaQXkxTHoT9tRPGuGkh07iHG7NDxJV667tAl9kmI0YnZqnvH6eJvWWUdPj1
smpoS1MPkR4J0AcZsR0mcunFYTwPAh4OPezlok0Ej+eWOp/ypUQON8ZRmRsNHyrnFlgJOK1Ufhi4
FsB5PH7Ws60/A5q9M7C6GluCReas0rOC+nrZ5vZbo/cgX6t0ajMuZ/L0kZmLrEeYkjYu8mqfEtag
j+cYu2mnSuqqVfALpNtOQ1pKTQZkjmvxI4DbxH4YESG326rPj82uFx6+Krou+gEgodJsWRhMbYq0
MWgPUjHUTSy0MRfpro66fP6/AMZGif8UJuGkOHJ3r1kZW0YNJk0ASO8QRqwrrtT2F+wAocqrId5D
0zvvM3fj1rgqKRT10lnjn4xpkbrboqhYm+8+f7GbNmFDaHcf3Q9L7u1lUsHLCWS/mDSC9v+cxSML
xLvSv2SqTIFMTJOqdruNpIhOiMPrO7vvR5iXMtTOAYK1vLOxFG3gt7UHfQ6y2CZQkCR2i61thStj
/fXd8oyuiKNkgXnOW4kkd0RY9Ea7HqcWhYsPjwNJpEV/iHTO7xhDRcwzCnlLjGeOV/qUCVMBqDYx
OcL5qOweNUEcQu0HDAcfI4K5cfI5pkSapxdulbx37PiY1I3hVSsJQQ+1Qy5F8xiPDNWwPXWQL/cg
JjQGYbWqIk6n21ByemaGjEBG9qL3Xt2OOXt8EtJfE/BUdtCsO66G4NKDzZI4tmMOZVjUnWB25JmX
RRZl8l7zmMqhac8UZweFDalZsEI9SGRZcso+G96CMq2WrPbStj7t7GEt9CJebvWBoaYQ7GPPNfRJ
+BihODmZTZuCCnGu3H6av0HDiuhIQusuj6vGiQh6rAogzNtOeuCl0GF4d2AvaIKay9QMqcmbcE/s
B3E+zAxrfzvJ9YNZitn1Z+x1NjXStGZ2INc3lejagQ+/O2RuYnuRJbek0eFfSYNby5ufhCzMkTOp
aqBrKrOHxmTMrr+6252wTyzJNePDaAI9eJsKzWBuWvch55xe5xg8MwiDg+dbaVp4ptFdeF3FcLET
QPIEs81AuoHsq1agaRsueUMlKIfBKb0QnECqf5OP5tfv0XTu6oEXBeF/x0m5qBzhoOHK7kFUb+es
N3pwW2eHys5OLMv2cMFnxYwqPAL5CKLe5pceGbft2aruCYUXiGwocDy89rhnsnHyMEVX5NYtTisZ
uu8xQAmUeI4eBOpDVNhX96fZZvE3B0BLGAaTbW7oqiUxiYHTKugEq5L7sMrXt40v5qxr8e2+dI23
zDp/7PkRlm1dwEqwK9Ik9GXsH6/tsLMdcnGrH+uEffxv3iI1h8YIY2rPEQE7lJgePiAE9dOD1u/r
lccA4j5jlAbRJPa8qO05oMQmgztIwadxr+Z6KYX4SOyJMxS+XgNCxEOReMi1IFPkqvoTtHFzzzdD
fQYPQFRBFsohhdeaUU7JNXAaM6Wk/gXQ2cEXQk622tOLIJxIvOf7iqEAPBcyNFluW7my34PGja0M
NqAOIsqRe/Y78tGMyPRd7Qcaj4+a5ZN+jKbu8neWdRtRVauq1pPfN1miI8U/EzWtWykmqjvLhseQ
r6FYWy4mMumakfumShflAQPEUaQvWpRhgzNnR/sniTV8QyoNcYcCpw8KxY0No/s2hCgKdUHr45fD
KH3qwIkAPOG0xo/dzZqYiOo7bcrPChViv7RhLEsCOD1Rto1YlnQEGRguxLfUfV6DBHP8VCZ+cI7e
C1ZVwBidu55/Y/a/jbZlVyFgwRjM+DhvcYC/4MQp9MeoOGu+v6ZNVgPyVp27y0a/jLf73IjMg/z3
kNP7NHCfeVei98igebum38xmceE8CcfXWt5+a/AEQnWPjdPeHu3qwZcWCeEZM2iCstaTewLmrxOs
NJ7nxhGGIqwCME3Xf59OfhVnIrPO3wm3ArJej+mKYJ3uS4/gyYhYQc090s9rQT0YLAWOB6VAj6Xb
hLPMMWPgQIAlfuvgtZRMlbXBqnU89iohp8R5c8TjFx4b2vjixkuFLil8M3hVwAzJae4rRkQdgffz
EyRtN6M6C+vigSYENFMJ0Ms3V+O+0yOoNoHaLvC6TaJInK8WH5uB3h3hJvw5jv/wCquX2GaXl5Bd
Yw//RmFBhZvMRsejhMy6ZB0eiGLkDNxc4X67UyYtdPyJqtAQCEpSVgx0+SLKJfiBCjZh4DnQNrTq
6M6Ue1A9zRl648LFSaym2CwysjAFvjmeihvkdtK5PzFdA9Q8uwzxBeVSjJ1R6epNCh0dw7AdZU/K
WRrKKGldI34Xw5aelFCed27phTdqGphKAAXIlnFRji4ow9QnK6MexET4bLvMXoCQdz9/12SCAzLt
J6sEoGHXSqEPN4Sw7g4gQco7i1UJ1aFUCLURfdBO376/1PP6i64fh0QM1k5XLFfK2FcUZ98s5KGg
zBi4ydmtboJGDdKP0TkT/9UtnLZ7ROzt0geRFnqsrQoiq7xEiuWRIHjsmqUT9gTKxG9JNwauLIKG
1//EHfLa2CLlGvziUna+xMkPngMY/IlT9jmPP5lRUtFqrR3E1neHGV84rCeM23WruIvXNe3w2Ox9
SwRba3UTpBJ4KQehaxBoywJs/+jd/Uq3LKi6w0yrxvAvjoGUJkgRts5W8u17DlFbQ7IV3t0q/Re8
SzOFIXLSHVzG2pKFa+TgfK4FqhCBI4rwZ2a2ELE+MlcY0UDu+brsF0091i4+ZqSU7ilWT9rU4BtM
TsEry0EQuJqY52MJRNtF1Rsdk6mZJT3Xs2rBTwDDd4eHjCx7Xs+tI0BEI6zC93NfNqF8udrGJruI
TwGibQAwABeH0eAj15f53XatQbqyW+sNoAU2zb4EiQmQY9taYwI9lrL2iivBtM+0OQBkJWqNA6BM
4Fk30yfrD2N3da4Oc03GN85Cfoo1qHIHtUsMKF/DMWHf7nfhpGzE19hK879hi5yPrI6o6CksZhkX
RWlrLmevkaGZDlrYzKOJM7XRsON5GkeKIa9PAvkK8GyLic4/jM4WrIWemd/FYgPT0hge0xeESm1W
u/ZuM9BGkFO5YhmDSaSCnGueMoOarhAUd/UmBw64ej3CD5XLt9Ey6+8ykGRg5J50D2crTLkUmkui
RfLQhrX4Q8wuuJcLQcQO3riUkkC+rrbTV2IJ3dZHnmmRFNVY8mv7TNV27bv0zHangk8IDTQmBldQ
b0M6I0Q8zA5WDzw/HEFPwzwUPZbUmPt0q8q3DDsBoepB9IJaIquYbL81FxafhGWUdur7rVVxpMRf
9WLYfMmjdoaIcmK4ol8CvfAg/DhTd9Iy2GeFNyVA7RTcr8N5LsbmQGvWQd62rwNjQ1WqKdNOeqso
Se1u4KZQsKzt69BneoMF+8ghP9tryLS3B1ZyWMQvS1aoJiuWHBQSGrEcuzE/wr/8Re5jRSgsGPxx
uN0Re8XrITBZfklSwGSXbW0YY47VdUeVcBmnn5tLBxqjS/zn0t23udc+guMW4N61a4VGrNtYTABB
lkPkgSvt8IkdqOKFLKuINupjPWM4LlRJ5DxJSGeNTde6Zxnn6lZTA0C6dtXlR/q0Dr7WHbnUi0wA
ak3gVHMN/EzydFyTwbILacIKOShY6RQFt+cjmR9Jy8wV6mFpQ04lCI4PQ5Ae7xbcqywOwnEDgIMG
FNxZOsZct4Aqixz6AHPznLeYL4qXimYb+hI9gl/S0nrGbHY7S6/wvENirwAIpf/dfRxlJtVAccGo
sEqoXTPSx2hwnhMYMYfOMb7R5dyOegMZlONJXtre67zTJ+vKhrjdxeH7PIdOz9c2gAheYel37Tl3
fuuULcLqmG8C/34chW8sDfwgeMIeQUJjhbAd+gssleo3JkFOIu1N8PbeaY1aaW9LtlyrkFqPH9X6
3YMDSZtBXPGTpmtQ1QwTkNHTqM2pmz6aF2W+nbh9L85uCczUzlz+v7e+yIqQuzqooXBl5JmxNPpU
ATtHGLe0a2YR+RGfta6p1cPZy8IdY1k10nhcykDErJf93EuLKbN05EjO0RdqLx0khtYFgRASC/kF
OQ4ssBMg1BS0XpshMOviEvkkmTB8R8EG8X1C5cv/vBqV6Kzxlsjpq/fpg1S6NC0cATXOLD4drFvF
30bp/C3otG+eiSM7hAC8ltCnBXO5etzNc7YPnJUPe8AFZiqYVWRNxdrnbs0MpG/3NEoaLDcmBp2k
gpjXdXnrGZBx5V/b3jngPGmMUy6cHs5C9C91aPvoap2DNJPU/aSgGhWFNUpiPliQOfFv+ZYyKi4n
d9YZJyvyux7jQR9v/R/oWm++2sGcMGvFE4ulF7bW9MV92cQm4hv9LEvgxW31pOcztwQH+AmnW/0K
eswgr7ZzI4k2utJXQriUCgJmAPDFz4u9psvEF55btW+D1KpsDNZYkNxyK5wUGqtrW2QoPpEsBVIx
ykYwiEC2wJ1Uu1odBWNnireDGp7Tx8KttCpo+WBz4hWXFz+V+1xQuEpBjxvwaDkdcWM684PurS97
wNTkITY9bz2rBw36UbCUPDyqVcjFXxXvEpJkytFUGapa/6mwn4HNbpTnAemvqQkh6ZKJ6GzWG0Gr
AvHCGY/s2oeePnNRmx5HsduKPJWjN35r40vKohUz96Hjtof9feCL/sY9w9n/57t2g0fDjnMqyLXi
FkRd4br30VJ8MVwM+fw8a2RJIVPpxwAfBGAupUqpAIoRoURXwbRMzg6bw8yf+raRDpZmtHb/LYkC
+GnoTriSuHBrEhrQehvF/qL98ON5F0fiPVKFk/r5ly/d7BEStuu/O2Y77pJQ8KNzAkUxcJJYEAFy
9LtFYOzHdQzgZbej40KBfzZF0/gG2pHd7TBaDw+wsEJSqTJ36qGYZI3jWd6Eky6az+0yMVqK6ubF
kFA5jK/uXa5+dE+o7EUio1ZOkRDqjePrmUWAceFCYFtoeK0dOa93pMq8fSq2YEnT7yMolsIJWB5h
IHLJxL43FRbRuHAkeG3yNdknaQKIJxXHpXEhcgyFjVPMJ5DMtguazTimiCdSE1vx/fD71t4UJWps
OGg2pjFkWjb6wRDIw/Tnf8XqpCMDBx9tN7HcI+CyBmQzzuP4DOJOtUpb7+B9TmNip5abTA/hf3xr
wl4YY0cnfaQzL/N6r4ZbsvAbrAGupkNsoc2C/CR4vNyvGO18aOiDtWwYAIMSTVwp1bA63VdTNmB7
rYs7QadR3jZbaQ52jiNkzBO/+y0MOJKqMB+/lKPa4hKzEw8/0dH+hzeTeo3qKiJ15GXDtYRGL4Pk
BY2l8kkyrsBkI7ErTvADUFiCBCPlmk8OvBKR1aUtg5hqz7SjsZckT6/dipoQaEvx2hQaeX15/WmL
D8cwHvvQ8hxLZEnLcLOjGCCfPhiYilo4iudtZmInq9HcDK76BQ7tqI2qX4Mc/UL0Lcam2P9GWVmz
xAQW8IkabpvcOhPfTo26Dtv+/OKv4Dk4JRbsGw1yxxHGxT9arL8UyLVfvaiijhjFpP+nLQVBgNY0
WuvNjJuMwhC1mSJKOfugRbv+bQljBPdRVtohQFlNsE+9UqpNLz+cB3pCDaAHYrnz2lOdmptWT9UE
NFvtYqY6y+uMYawKMDy75PFqmZmGTGEpZgoK72f6wm777LurVZnOWoaPt8k4sYwABB6Z/55uEzKg
NAjLXIPVM/F4NjBSQD66ZqZdJu2KRr7Ek5arS3w/OfgTQK3ts7iFKkseMnmKOYzNpUstjMCtZ/m/
ERZ/vfcdLeAVdwNHOCK5PDWaePDIRjdMnkvTCZiEkU9Jhq7f6v6399vM6OziYZ3kwcACARQ5L9iL
WxeblYoyI74ng/tbAXncQAzKLEFr5Ci0Rf/1Wg9WIkWktmVt5RpDi7VPsN23YClPAoG1s1fc5pIl
DW8W9OAsbNdAuDIxKzIl37NRsF2vwAizY//q15mFD3LmVrhl3QMKScLHX/RLZLTGF2g7EjLHk3TF
cd/zAjXfKgtQ14RHf/B7/xUvIuYheZIptKhofp8PcqtKpGBRcuaOpAF/NvKHmpfFKicWGo7c37R7
86SCfS4VYqxn5O93cin3V9j9s+QAioded5i3g98xKunobqmoKpT4a4QDiiCWtSR0rnlbRsQHT3T4
5aihFm+82c4FHXXzODfSZ1u9OgFB+GFyshjahHYNupbXpepLmTHfxNDUNtzOTY3jJBrU2cvAt/7O
kgtUH7GGDmbLB1P3WY/C7DbWN+t/s7uv6KwJYzPvgPSSyZBvDLkrOb050CTMXop8Gpie8gTSC7wh
6jj7hStKdPDyGW+EH+fgQyR5Wjaug1kK7+4XAgjfuO27bI2wnNmxMJ6tw09gmSpRZFyGpaw92xTA
0mo+7QMtx0u9bGt9OywBrLJM8ZgEWcs6tRzwezidcOmWJaZCN19YhQz5JF9wHNhz7xOmI1CjTjg8
/TszFKNyqp4jEu3pv3h9dmyFTTz3wX/hxqyGDeKN1pr9zl51rZnUHzo81umwrEX2hCx3JW2lr/9b
FL0aWpRKaV9FGg2lrRDtDRWH9R8+uzcnunHohqQE8/vdUj0qTj1OpaX9LxsDLDhf5GbRoUizAvtq
U44E+m/ZL5zJFKhJTmeCHxX2Fj6MYHMc8M7/UC5mOVf/A4V6HUvvvgjY7n6dnUgo4KYmDMnmnohR
MBeSBD6qTestsmXnneTAjB+jkP/rojuZZzf7cp8rGqBXkNWMMW7jfcmtzQCUzMVJgx+OY3YEIWhH
pz3KNO1Zg0QPbUCqHYF4XBIAGn7eM2NFyQPIGmGrfLlcKgOp0krbf9QMEKSR8+vyId3EUjBuke9I
3QggsVvvLeaiOm4hWsay5WcmyF8HyCGRevEBK7XgKFJDW9iywsAxwcD5Sj5m7ImiSU8x9+pWINh+
DWoe1/AaHVCViAvGbwWvaug/vnbNjHmAmnSvBS3uTsD2nP/D4Xk/wUXkM29B6mhjK5/WZsoUrrK4
ZJpPhDdUrqUXguLyfAunwU6VxhmsH3bhQLd6Y/iJ7bCVe/PgYDTGCjUPpawrRY4q7ENKbvO5/WAE
9GPow0JGLbmK8PW2OAgOsBFS6+zdHdVB6Y4MopWLNjZ3SwdZmVF40kcsfzstGy0i68+SgQtkivaG
74XRN9ubsNVJ18juuyh9AgVWMj1ciGAAQxxairvc07SI+5w+equmR0jF2JiPzOnD8WkjjzITwSUc
6VkAr1w/DrZ9BFGAYWYMzWBqGQhdWz8QBBTkkX6pp3dTmO+C3q2xkvqOVdvAcqXJE9TUMLinyetz
0NGf0FvoPIK/cj+BH+17mUr6wmfkeW7QJg9CsgyWxX1ejVqb1xyw23WZDJg1XSN4Y+vIM27MApDn
6WzzekxbCCXurBeNXWCr2xErQKkhxgWIfZM3okq2GtRLzeal0CPLLw2OSceEiQQwY++McaMcOcLr
k3tPC5+iOPOLOPg1rGZiIub/+UJcyYVE0oLvhZHT7Uc7Hr95aDtnO00GDgbSiz3ydwCO25Y+r5SI
2HL9kUDg0GWda6p0R+5tRlTuIeY0jfR1rc5HzQY8feDaNUCeWu+Xi1PFqh0tQhZvI61dfHDds4Ua
X9bm1bi///UiITR5jQxQzp9aIS/OykJngT/xkBZGd0aDmGTBaij4yc0+gRhD7AVavzRfJ/rAtyz2
8cvQkOTVpsQZjfre3Gfz4qHur4k0PrsNASATb+HCqEclYCAyRrI1iJkV/JMNB6GX4T+BpOGrgp4z
inTq65BAHpFTSRZs6EAadKy/t9ZGe9siDvR68qOE0bHSldXFZW+WNEzXP+5I2R9Az8pRALxwQ0Ux
AWl8osgk/bt2FjpHNr7mRVjQjIiPVYWYxKYdXRPXPi4eYYn5z5hPcBU4+YWmtaO/wjY2dfBwFnIf
0MSMKZRR24Rbad1S0sS2b8bmjrDz4JTQySLhPaJGpJd7L0O9RvvZ/HD8wY4jHxFU23V58m2Olegz
sFgZZ1+kw/8rkzUBFOeqIJplfojOS7GBKKVsQ60SY/Yjw+SeESwFu2xt8dmC1cHpmi+eaHjC++2f
sffVB8/+WwUU6gABSoYJTXBRGBn6dofYsHX36HmC5U01X7+Pvbfg1KuH1SPWg5ni0X7ZZoA0Cs7M
GTF+Ljod5VIz9ugMZLciUIfXdpaxB8pRQjSUwpd6Ubd15spUguON+7WJ00s7UQ/A/5guaR2+Q3fJ
74GEbUgTLAlLCa8tsNqI9LQpq37BAdnf/1sw1itJQqbH74URcRtVH1+U/ziloPgyARQ+/xE0+evI
RWLCenSwrZiG/fwZt8CariX7LPPURz2F+NvvWpkB1E2yKQBulnKU9fEnwlhFnXB6Z6ezsUfasgpV
0+5m9z3jlFHQj6rpzYxa8jJFmQrcIkN3c0F90svEnpDeu8kiwoxAZj0CXU+aGLrwvDAmHnmphNNH
FywAKctdCB0dsIsZ6p+W78K+69kBAAEOB7g2MkMY3eCKdI+3X1tap9Fnkzqar79xoKloHXMMonS/
9nesnRqct0OQPfcxcnqbJg87OaoUGPVGBIYs+Iz9chOLERAZqvJ3k6/yhKLIwv9z9BtURW+KyJ+7
NJifGBTkf8M6v/qtaauKTCsROYDbPyAKkZyYxi7fu3MJOXkPoqpxwCtvt2HK96Abp/X5bynykvuA
VWr6lORcJqzpOaTnkLdjsCo/WyTrTzILbDERVlpJjf7eoC6OzKg0oy6HkJfYq6JNE0Ql7AiFsWeT
+/9eDwMm6GotyJMJ53RQcE7tFTJ30H3Koe0R0mto+KgXXBFquRYVQwXS8bWlN9ugAS4tJyjC6D/W
gOzwfXNGDWdK6xySeCakrmC5uw0flkLEueRX3KxgWI3IdMt/aPag1wJG5HLFwCBXz6N1JNTZMPos
DDEnMB/kjij7I/DrN8nv9H/uzg11uy0znHa87v92/2DYCLzSdlPF0UtUjTjW0bksqsKOvnI21O0I
9eBWUim8QVGpkk4fZshTz8xi0+c5KjK+brhiFFhLjBYipbG5Y9bDQdx5Zd9ENTBKVffrbM3Sq2bH
zWkix4M3vc4s9AkOKeyYRC56PGtaS8zZfsvUPXcBFwCmF1J2hmdjyhImk3ei9VnhKdbNIEE44iIw
VZXewVuPIeogsaP73M88wnE/tpgm39qOGo6NsMppsOx/2T3PqoBBpj508saMlE33/C5/1w7To11y
lNAJDeJcsRtBA/PWvMpOMVacQgGUkEDN3vY26jsP9LetXDPnHWKTBvdNAq/U2D3jOyapA+LVQcU1
19vGlJvEIzUFXi734FwTfJAQrkMFUb8TCOG7NSJ76ilXOHE8psfdrmcjJU2w8uXiioscpIFwZMSG
blFvKsjaJNyc5wlY8yNU3T+Kdi/iCgZQPm6XJO6tc6fTollYf7RAvP9MvW61XUanWBCjxnZIb2n5
fxZjJbq9xX6URlTfYM2vsOZEtpmi+zESpsRDSlni92JoSZkjg1e+3zY/7eF4wcvxyu+Y92BRwzc/
6lzunJ5nMrzbI84oTxZb2x/zm1wqGp1bUD86r5quzr9PNwAiDj1MMWxo3+Hhzv/SbvinwjKuXXgo
aOxgjIntUmKJwDu/OBO2hR/WgFz/ZO8GcNLYnVNbqepZRIBd6PDTUn9i5eKxPyMq95owFUxb6gyi
wCi449bAgldOq7vXTI/nbZfIm5yq3BbTsleJso+5CICR3QGxETH+EybA9HK26Ql7TAnRjXxyivjK
urtUjU6Kedfy1tuj4L507vKYsmCjPsjU7G/TXQxSWJxrG7X8lZT4CNOgEIpZnEa4QpJDthbcY5xl
RdzpWMzUEB48SJGWiYjWGZTunVGcZ4Gdmv7p01IwB2kbrMfuMlZ7vetw+eoTbKbGSlnsDLsw7GkB
Vt9RS5+bFfVHF9bDlfhgNB87xlTpUURGEGUOJWzjGr29lMIGkeJn8efFsNHZqpVGmE62By+fhcrk
Wv/XA0A81mKMEzAgBGHSwroleBrMMjeV0OUQxXg+WgZxur53FelTfqlAnn3hIXnce0hd2jhupPpK
1h5sg31+0kUvXNOCww9RaK3wBuM2QKFg2ZnVetaoweoDKdbpmQV0MUJiPOEFypDfysC0na1Sw+bU
QlH/tgCt/mOFcFZcTK+UjEPjKsg4Zwhx7vPrC6qn+JxBq8h51eb74xnHppqHj92q7nqZCgTQ3Y43
We4LqY7roAPQykwNe05Mc1lFZRWlCHOFGsYQRYY2cNr14/3E04swN4Y7o5Yp02iOu2ZVK7ujisrv
uAVfrhygDr16glVSGCunOWJ2qZqMLnIpJq1k1OfzpatbtwwjD2i2Ndg/GMyWlTP7GG/hgCt0zwy9
l6jp4ectSKEFR4lMhQExUQM7sMw366mBgK/IXRG2silRd6J2qReEKZqAuHsPPFj2FQjdeln9GjC6
UK88cPT/RRRp7mE23TeSm++g3yz9TmKxI22Ww/ipaqJdMt9vW997TlyLyzig7g+0lJrvNvc0qj1A
fNK/MsGKYNBhyz7cZ/SR2K6fQnzxLvtBINWv+7GgHEBGCNh44y/xfYFBg+vduD9UC3MkoV2Ec7ud
cB9l2tgQjQ2guwOw8BRGkUAkS/1dJeZK5u392/+dI8tF9HCPVO5NMwNT7UTlyiqAUAzDlkcwRC58
4dXoXAAP7dN2RFJ1fCxkEk15mm1ptcLICtoxPqxBOlUWfCD6ls6atE1qoXSccC31YfYAh69/9VBj
7sT/kOLC5+e6yN+I2fuHGglcQrUVxhG/CE/sb4bSvSXX+hX8ZWm+tOWaL9zwtW/gB+NcCzJ1EhDw
iNJq9kx+09lx7rDzJJ5Gu6/vj6XAI+GBB3JIqdX9g0wR7ALxviIFIDcj1zD1BKMKb4hfjtCTLj12
eIUepA91KW11dvnF7RiQQOF9BPjEaGyh2RZz9KPTlPbJf0rqFsgJxFR94B7BAXR9mNpTtTxaAP61
nSF6UE9cLbn7yTFqbMBifNXmxtry5/TsHJHFs/d+yiH/e2t4AI5triqFlCLpbG1Oi7gieXJIR+Gk
iQ8IhbxeiQB32fiB8RYhOLf/57jbrkpg5+CFJV+P7M8oYtm4//PmPoRf3IgZ/AonNWn0w1FY9jfS
aNyx2LfBTV9E9/aIw0Ew4BASFvY09nuhoe7X3/NyPYG2jpExlpg8Xcehn2PHKZXRj5E4NHlcevnk
W6ltaKNS+lkIxhC/9KqDfKXf8XOBaxCSmg4Ajl5rmQ1vHSDniNhzlX6q8v/QpikExsV2lPkavHAg
r5yTwjBiKLfYSvLN5y8+YpS6kz1WUpSmMquUbNX8WrMBgiPiN3oc1cCopLuJYNW4FDZCs5INm5Yv
CUeuZY2Wb6j8+2DBsRw5yPOvmduKn6LaQrx6pwtRbq8NCfYuRioQO0e8qJwcj+B4WhFJ3C79i5A6
Cpfs4ZMkPwbap4SwQV7rOlVOImHlOp+gCfpBThLgS4DU9+VIfr+BWL2D141lSdV6mKn9mx8VtfIh
WYWUO7mx4b7k6LOu2CepNpndbfFglHvQuiN6wLD58jCXvBUBLf59U+ne89/lZ59ScFeqtGbG90s2
bQ2HVRDzaPG/WHC+Q3WUdVhxDOsRQZKuB0Y0BwI6ryviiulkX4aO9JKt3AERb8TxsjK9VF6opZXs
CvVsMjx/hFP7/xtBHyZdLPVsBhRTKzVmMTJX7nE35vDDjJluNajAZnjHReQoUEEqq6AsqN0vhI/d
9HhhhGQ2hLOskv/0HS8v4P8/IYGM8mfin5HipkWOQS2VH9g73VK0TNyFs3y/pSanHF1Rgcrzuk61
8fdldKs2nr8mlJEm3JyKHZKwu+rICKUD75sUunJHmFRI38f7NdsedCE/sMHNSRRcBXu9J4SX9SMz
PqP5yO/QaH97OFJEaSQGFW33fc2YOBaXgC6QAfMX3b9+MGuQaw0CJt6cRavI8QhJbYHDj5iBGYw0
BOx4BZos19x6bEyTHRn6C7HB8D1xHaJuIw6kOBMwsSgD14NNhedD01qrqdcLOHUptPXo9afCcFBm
1VzGBMXZdrJx+w4X0BM4hgiUhQedT0f/VvSZpFFCuz/hzQzrKvWPMBIrk2L4zJp2G/9OPhzoye5M
TDYQXwvCa21hwEH7pP41AK4uDaRg/5C3EDLseIifV82zolPVe65Tk8d/G/YbuMj6GSuLYwPwd3m8
7P/xZv1X6auaiCsiH8NSCNpfOVWq6wSM4ZQU4x2YODEgo83h5xxe65hAmyRjnncZlCuOY0JhN3qA
fZyA+pMDK0eh2liNucIQGZhcvJhw9l4AY/5nph3avenNk+xciI3ifsKFR30PS5/46FH5DEvSGx5f
6AUDSf/iCEK6pF8bOulKmgwYRto/7x43QyTkma8rxNn9GT2vnoqTYvcx4TPovUjQJzgKNjIQfgnK
E+MUxwz/L8Y13UI6lPmjN0pvsRh2hbd6BbtgaP1qznPZq8ob+RBHGdpDstkxntKlpAo0DD3lzS7x
h5fTkbcBu1frUOM85RzOUQQjJj0sJkUMGduQ9Mrf9aGeyE1wNKswGuS8hLh3TFSY1+udB2IG9jO7
nXQX8QsfgIE7rXAiYaRoSnZiUvR3eDlt6HCat+6Nt1JPz6Q50xcWHE09rVpHstEoOyc7ju1DWX2z
LlFvHvP1UbLaYvqGelWZadyO4RikGoY9DRH0uFgCUGdVd7Z2j+0RFkhcR2e3QMB4Srp/IUSyl0Bq
DkAyYRUiyJ1PVpDgKTZs/iyGP+h5GxNwYfak2L1i6DdsBMxGykmLgunU5QtirMhtU4BMxBLwowv6
XKZA+I3hsCeRDUUOTK3Aisvd6QSR0mW44RYNFGucS3JrTLG7se7X8an/Jqd2USflwGhNGb1G+8Ue
yuo1JWnrZbv4eGrwusrYLOpRjpLBIOEsZJAjku42BMBX29TVqbHk42Yj8Y/f3XFgM/DHv5LBwBWR
7gqFqPA0eUaD8F3LXgRd49zvvkksYzXNOebcuOxhegXWcso0YsBxlLsQSAQvNKeZ78rYBDUHYQQ5
61CM7viMijKlc2+Q681s4BMbdhNrRwrpC254zVudJ4XQqQ/9y1ytSbBQos5INlTzVudfp0whil5z
dJzOXjCFT32OXfGNl6ruv2AZgGM0jaBnm+cFfI8glXl1gzbiJQU6uD+YfFD80aZwEazpaMu09ox8
SBsPqB+giHp0jwBgdo6sZcckVRz/rHmxVp89kteIkA21fd+SX2J9J/ZvJMsD9zqLuiRJTuEBS/aF
9L3W01j2eJ/Qd8fjT4+51Y0vLW11wljKmGIkCgmaQjiptIPMIrgMtOo1R8qWm0rkGZuyvsktu3vL
FmxvMUF5zYl2/dcQ2psZye358z1xCIh6dnKfg60XQ5RbtvI+Ux6mpMdO7gN1FVj0ivpWNL+Sax0M
l0DOmfEyYTdIln/QV7Y1/AK+6oMtwarGRvKkm1IH70FLkziWsA3Syd5GbgQQtDrjGt8+bmn3BiTv
dr4IQ4lEZghs3YEbRCQ6wku5GIbWk6PkYuEyrSxyj2tAoB1LBhoC8c0IEmZZCSjfVgpHXlnTFywm
KeDXLE54yBafPa3+wxOg6U0KzT08Im79cqUWrSowJZ2ONpQs1Z1jfYWqSMCobHqn1z5OaBarz8G3
m0KcAgqFs0kiWd7Vz9TKtYmCka2elfwmi3nebQ9bX7Q1unnp/HjtYosLGJUDm7mC405RFvYdVWUG
23BZOfz6Sx9Ee7RqfwKXCPS9wOcmu4Lfv5a3y42AxsBFfWTs43H68LJkTmC+4QqamI2iyZPgN5Rx
5UT5gXWZ8zqlCnLudQ7aCXtm5WgWjCSduhNX/btOQQoDZnB2gf2Ot/Yvnkx7U1qSzS6bD/yXEVQx
J3IKM5bbpO2bILnnnhAA5jSahlyY7Jc1Tsf97/YJngJz9LzDz9tngbsOfl4PBgPsAZ9Epw3ImHDC
QbiooTuJ3mHuDZKuNaY+ZQt693jyLsXS49GKb9cRJXoPC+p/c8cgk3Wyy0gzmfd7K1ShAtd/oUXm
nOZyGLy+2/aBfSzqNwwQTTHq5ZLPCFEbpmAdiPxaX27pWquVq1E6+5KbQ+VzHJrfxdn10j7sHLDC
04VDHADAaAMN/dbSlKM/e4oBaYLHtKwUNvdQNzPkFNK7dBleXOLetcj57ajH3jDjPe77YCavfbFx
qZyQ1fv9aUy/xNunGX1ZaLaE47oy5iBNsucBf6dVMR5TisA6Cnqb7N/GIlvE+qEOa0EN4E9kyM5P
oe1BH3AtjpT1Xaqdm92ZvfWJIeH+WhV+NLcILqNV8X0ZRQ/XQX3IjbFhTL5QO45r0A1OlECSc8H5
IONW5IIaPhCsA60yhR7YCI8b+szkltOGdg0hjpZz8dxHIzmqserr2Xucpyl8PkLYNdISxKfhjm8R
bFLJnrsp9ib6j9c0PyKJfpa3bQ2PzDnW6Ku3qPyuN+APhY/W8LP2K14jcFbD5I/fY7vJzGWHygcp
D/rdx75TWk/TzfNzDYmi9zo3K8eCaovorZM5NlksiQeDW2ePc9LmLKgenMId0foJy3FhsVeisjwG
7oH/nkth6yn1qBkdKFZt/f4di9qS7R41fCeRL80/cxjzXm5GZiX8898FU73hxJ94A3XG/yJFrFvD
7IMrka6Qeb5b/K1HTIaEmrMkZZ3Ho4YSsCX3tTWaONFPgLKJ6PYefOcCRTLuPnEOcPqb3BnhI+FP
WoOM9VohabcQugE9nhaQ2qTWr1eO6/ZZo8wKS/G3ug1LTZIUcMufK3OCbDFbhWie8W4C8w66XkqY
LFuj4T/CaZR3Fp8cSvXkMHntvKH9SAU76QcDpxPJj+EJ/WwL/YXJ6SKjN+XP1ZIF8nQSRucCYh4O
gpozKHBSspoLRM5JJm9nteAkOKekwY8Nix8qlnDPC+bAXgTgwVcVtASJa+GNhNfZxCoG7y7Hl1Bk
hg2hBa2Pof5e3CEdhw1foCjmhNT9Y3EQkfMV+T2nGvg79eVpZk+lR+ZQCR/Hd7NROS2dZrSFWOp9
tSI+ktrCqg07Eue6/cYswuyKEvj/XefdzCZQj+evwsof5mWqxF6+fxXzuLChBQFf14elPcpU51gB
bk7PCMrHYVt2ZnM0Ba1uUzlBJXweWoPQp8auz5CeZPLvVggq+hpSh8dHmBrw0++LMPESauJLRqE4
cl8I8cCWpyHSwM/vut0fIdxBlDyWJuMu0T24vM3Vedv/7L+9g2oKOMrUMwOb+p6mD+7Dk0i7bAUd
+HIouDgGvcf+J9RRAn8s5ttt8ayGPALPguCgNt2eGJE31T7vM/RDIHrFbo+U15fVEEwDRMOGmhco
fosiQXyTDja83gJQq153AHj/NgwtuT1/X03cG9t0nI+3yCh7AVf7nxyb3/+/r71l8fshpA7gNX1S
p7BLkVX5nJNfwayI6o/vIO0YYtSejXLarB9D470OmLk4UOjoZwT1ZVxy0ao9H6k7DAO4bnR6ydy8
rHtQ0BFL6+lxeyz+8IAfXCkqQLbTngiRAeAUwFCaPFHtiJgiMNhcxvi3yy+2GbNTDBY0pgR2GPS2
vgoBI6pAtIpKMbLeJ61djhFgRRgCBGp41KmZ73X0VB8P7BItMSFHOoH43bAxYTBjBUs4fIiK2LA+
pjnt/nyznd/t5cZVPsDmL1gQTmzRtuztBI4aNKtLXo30eT6Ch46FP7B5PWIhe8TJP3Ey5IKjbH4K
p59ID54LGSYIAmyle5jVfqNGdPmpaeLnLbKwg5rh9vqbOgOWUEzM1CnKE80f+E9QY9pP4tBMHtiy
4zjSQJ+w6Bjm6yO/0U46tLDzQrZcPdLCLMQekYSrP52l7TWi71v8FJfw/jYJgO8ijODbtSkBiecO
ryFMhbyataLJSBYt24JXgXALXuTPTCIgPi/MUD8ni/sdLgRT53qlEr6LWf7UF2jsSQ8hROLrSXx2
BwOgMXCXUG4TdhG8lUqsEMMAjeChLQh2ak/txtd7ZLTOdfKojwBIBdu5535naXzSzjXppRO+/VGu
83woZR2MlXp2/FTP+ozI0khtxzIGEW/dHvpxZXecFw1GMx7eUBBa7FVNbJuKZ/mqYYktXHttRDfu
TwpLoig3ffE6DucSfEkU4HHbcgHR8UZ4A12fPWWOiHxlk84TV97ZVCjP2akggb+mYhIVOdKt7F1a
S5uo8+HFU8KhhTvtEizo8QlX9uzB1I/LPIVEISuaG2sW3mU5DmXnsSoP3IxJHysZnv4chAVVVU9T
HUxCWbLlaSyRlYC7ucEb+mDh3oPEla+2d+k4+/byeo9U5RUe0KWqkz7PBMIAW2A1UN92wuExeyte
SWXpq9dGmZJtKFK1XeyYE0bHwBqwcltfwPz8IFG0be/SapV9ItItaTDRbEzI6+1JHeucI2ZhxeQ2
BkyWOTPWJdeyZmWnIlj2veL4tlWpCkz4ISLINPJlD2AJQZ71qPW5aGnQSAlP95RZBhENT4KWu0jl
YS8Zhy7c7gQu8AOc7YPS0I3N8bY0Wz46L/tPfSnahcDF9JxLFlJ/8maq6kVBYcIK5/RrrksqJYMb
92KAsFT3DG1h2lJV7nKV/BerEDThIaaJAwh7PcUaLayD0Z0lYL5hOKMfYZ+6SzTS2qu3/GEnaMLy
JgE0ttyHiQ2AjfwPbDuad/HJsZWcrN54FDeeyHAqaDZIHsZFCYPzFq+AO0CTuphuon+7jaA0kCou
ZJ0LmhFJuPQ+bUthUbJYT0CWZq8yHkssghNLvaxsxuK6XxAOhTVXtx3XuznF3sjmpIfdjC+G7t6H
cbJbAIQWL4QaxpIFeobrqwcu2GW6t+RNufquk+g2D8t8ftY8AWDv5DIW2ZtdE7mfi2ycfOLtowgX
La7d1wfJiLzKEINBXPI8u5eZcFTo072yUPBa1CGDzEX2qVID1Gs/SuC4xIbhsUXE0V0vS+5h8Vol
ecrgZ6HgPRbs66npp9h+Y0p+48GjQmFEkYCctMPpXHH5BNUlBSr0G7g05ZvthjWo4we1jSZwMINJ
NFdzKdKDAmwRrEu2+7xCtsAhDd5wyt1bLuOPpLII3E97V6VjOWHeCp5JuCtQBV8SeGxp/tbXwEkE
zv3KaCdgk1ehE2P4gSCn+VBYZvx1dImVVRs3szDqoJ1TCO+i8G8ZNE+nJzkhOmYmXjXMLFlFYtgE
2BRrXIUh8aFKtIrInqF60HVSM0Mhre36FnLBv5/F2IFE4XS1j4iPtogJs0+hukE8dAQQHXNLoWCS
EEgTo+AodalqC23FH+N5umsMPrmIxchVTUeIqWv01iwRzh+FPLgOF3aw1SL+xM1VZxdi7cVbcgI0
/awHSo3S9puUAfK8Gy09d2GfjLq85Qs9xOgbz9jxcSxukCbKMxFYLFRJOaTbfefKEFZCXNcuqyIx
cJzVJj1t82E10Z0NEfYzdjv1Em+PvSjvmzMaMCnpUfWOTrQ0YTMOdZMFuqwhjjgytz7KjNetIZbF
lPRJXCHOJv7M8rJbcwq6XZMrgTctGqBlox5CDr0WVZe+B8qBvW6eaI3HPpLOsFa7CdPc+CgG6Ls/
AUonDAYOmnDoJOHu45sJ9A1+eZlqvIWmVjTeg+ThItX8ZA650xNZqNB1hp7mVG8b4mdV9tdbIaDX
J3QK0LTxo6yter+h+HwwzwinOkfDOVMbjH0jWG96EhcHBK1yWum3K8FuVfXgz3Dflqz1vdlCwIcP
/CYek3Q62WkxfkGTdal/n8bpuq0c+uzwHZu6Zu3hfoJGpqVzscMcTx4BdhaJ8R+QFak3OoP5K+Qy
a7ifD+NgkrRTT1KVYE4QgLWyRxw7tXTL+9fqm5MnvU9ei573vdKBcFbL8I4LAiycl2dcZiWUHl9d
sw1AvCdiGYu9klQZLim0SVQJgShIexMh5jpIU7U82U+p80+iCz9fne3A9TVaS2g8Xg0BRSr552ex
HmOmBT6VfWG9JoCw2FG9xQZ5VcqO9WUMSmMS4i3U2CSw5qg7djDKLsDDR5bU4eKl7tTbBlW32oD/
/8ilMhn/Df9JxTIZb0nTnZv0Dx48ZVOS31F9npoNW7Q0OW+btxrX0ekpFBOa0ZurXhIflV+Nwo21
I1Eg54TnIEv/sTJIzda+dZHY6ePNJL8MRAy4PCLy4w5kZuyjCVvfnwZosLf/ibmv6VH/3D/3gwTQ
BAx5xLwcxe7sctkCMEpw37udFJxwkE+wdCVGBSaPugahfmd6lauk6Hes88FVzyFtBb3tThNOHZG3
55B6Gzd8DKAvsbgLz/SsmKy4S2rP0qFMcHSvi4Hi3zldc7DEoVuV0aUQiS2E+bC3IFfbzxE/63hT
/fHbnAy/vAVOne1BxybXAFP5WTLPT85l6JyUGBX1L/ecly8zsRsaTHRWSQACFnDpbpO4/vUHYGju
0d5FAKyXqS7cJDCjLKKkWZiK0SV2JlCxhAYcZ8NVQmjg6Ri7A5W28GQe547F6CI145KRngxEqbTd
h4xbHQQb0ZDmJWeKXUDb0nRVlI7y7oH/DsrGB33MVgp54x8ip9a2+/pq0ns4U0d/TTrFH2VOf4eD
0giHwde6bh25MF+WkYS+JyKGpOQzlWJNxUkR+MZqDEuVY/vZhpNeUMfD+jAbZSJ/paWHeb6n+uHP
XCRrh481M8Vsa9l05RB8AM6usQt+EIoJ5saWJqEFkyAoWAA65GTAbTiu+/vQXsPGwR3KmzYBBaH4
qNcJ8aQnrOwrRxh2VqkDxxZwlV7I+br75paYdOXOEtqPCIqRs+3zzzCy8Z6KyVgHxdBeUxcmiGZU
7Frv7SwKhB25xJzfo8X3r4fofssyrqXOTXZAhicyyoffPuxR6AfA5xWWsbbIo4z2iLp/dGG19MPZ
Iwuidiv3JUbzUWAfTYKcYYCzuVaVgevCuNWMFX8Z1fEG8sODJSjpPl5KmxLwhmxAiq6I/lbsw/fA
XkHIoFlFyaeBk9fjDFm638U40JGAJ+Guf4kYyfNHfC+2QM2g/qkAiGbtFIrk41xYOjlMQq92Prz+
KTl2XLfvGvyxu61peAafoAKvFR2g7TQvgXjINaJhDot6vy9QrCS1x3uHqMw8YgFDYqIYXo9h/SHM
zZSrNPe80rnGhWipdlXuk47g647ak1RZsy8nS7gknb2gG8GeVPfRyj/UgjBkDOeEiyTkiKfdUxg8
vNej3xtYVzfImSI/T+jzBlygYjWtbPWclTeuq7U22ummd1Y1yJQ3qMjRjkHrjph52okAm39vaeds
kqh8FL16DiIpaHc23ABxSHC8LN0BIrgMGULhoIH6bBhoDT8TqWTfklwClsQX4zX2h2ohId67yFSP
XKsZjLm1Ilku+8be3GINRHA0wqbnjjgs8QJgDR7Zk8HPmzFJfUc7rvIO7ShFklFbQUpQoRTcdRC4
bSWpqnmQ6ZMoN28Lzulb0DWPkK75g1Sk2mi7k59HV0rQ1ScNN3WatcwbtuhFWAr3oXG401yFO8sC
PBA71KY9SqF+ZwpviczHZaVRy/1fm8q+irEbkladYxlYuVLO67YTaVNFj139EQlm8LuB+tjIJ/0p
HIGsbqNNzQnRoGA72GqlaTb46wogDNqN7yPRQHBkyw2mWpxzVYe0mPo0f4MxDGCLLeCbTaken+CK
Z3NzhLt1s0EPbKox9vKWNPOXNWycHZDBGcmCxxgFdqz2ZIcY6blG2rIpX/9zepyZMyi5ROMUlWaE
Y5SnEhlooW7W6P/ullIPQ2zI7URt2loNQfpmAmc3EVHrqKtZwQvsPt+nZywAlFHCe4sfipzyfZz4
3QyUbx+I2yKCl4y5L3yd5K1FoiywBw5tEksXnfAjOWsXCDuL3FArfcyYTxEbTgqPrnnxJnm99FcN
w/mVu0HcbtQxvjbfBO7xnxKY+//WbJrDsIJ7SOt0D+Y2ZWDb1Bpy9mp3r8UPmhRPEOCPMerihoDu
hoRJ/56oDWfiO0r1Y9bNN4L+aFI4cVqM1CLXMSRhYYGRvX734Iln+JMFquPVvFBTS8oSvicwxy4q
bBiM7GBFgIbqdw4Cxwr5x2b5ZVCiGkcmaPPH7Uo5BCcBCNbgKG+eHsiWreoBzoDx3fQ3wT7u1xUQ
o4pEBo6g1uGKrnWAzMRvXESTUf3795fIc+Sk4X23qMWBJluzXf+OfC7fL4hXWwuXX6hoyrpeIoUs
hDh4xcL29OWA75udTqWx06zK2KmjMi/5vusZdAHE+xCgLwOtS7rzayt2UxX+IKc5Sm/j81J+ZxHD
IVpJJp6o0iDo1b4emhepjQwb9FR23cs5fsnOGvvPC/jODBhcCYKqEumyiC7fBpFTKZSCbhumtgGs
l2ppDBCdpCo8eNcPE7975cVczR/oupED4wNQ+Hqccu+SzvK1N4mhSOcaBy7oFE8isxAG1YpIZAgF
9gPUo2hVXrIqj7AnEhKVsxpZXA6F0pU2ZB3a08USZGSbw5eQ3DnQFKL0XDIoqgf6bCmgDSZtaau4
0Ug6tSWL9rSBXs9PLtlKw01+vQb0a0YJ2jUAG7LFds9K0BMvd4LFWq6J4+ZheSHkV4E5GHUmLIyf
AAXwnxIiharOHq3xo/an6pVnVrTYiuN3z7CX9/2z1GR/haAxUU/hQmeJCx7K0GujAKdD98VYPzIt
GeiqzXYQNuj+niZgFib2qCTHSlZmsjrSx3jLRB0hhwm3HCkNZwvCc153ZMis+3VM2GlaKTr+fzri
23/LvdHyice7aLh2BwgT0XX/lGJRV9x9p9PIe0bbgvhw7dRRtGcz9nvdNRtTUsn49vgR5ogd9Xm/
9Y6WuzPoOPx/OO6pVg1wuvpfyo1DJlA3YFEK2WmyKzGu0tsXuf7oqBO2UBUi7FKIndU5SRfOfgLv
rG//9FSZshi/lhGUa5tpqRU3ShNNUcQ13YP6b06/a7OpLoV/U4lp32lljhCrcBIusmGG1m4/Qw/F
XXM5pIkslXNu+PC8myiyKy54b//DfSh3orz6mHT5DM2ERCEs6jebZxnx3tqSC5D9daesng55mMfp
adIZErN8fLmS4+y5PF9WR7Q0kPVyJMZlRV+f3yp84XgkEtyT0W1XkA4xof43ildFmxgt5nCpX4WF
BJo8CtwHgrlk7gWoDxHzzH+D8Yzt9jpuwKOrBLOazaAfEyOozmY/PNEsq3oRxjDU4ia/erImDTGk
CZzz517k8LjDrbGcbM1c6Rc/t4QfWLeSJHKwNIFWEr5Q8S51Mp5z90MmBh0NXHJhIdli0kcYja51
HEu6FVwSh8RO4Zn6dwfUdzSZIygZuJqdYvvyANM1jLJ5EACefMY1PoDDUEsGagpzxqD/Qk2WK8s4
NKHJDbTeA2Adik+sNDYbV6daKKRUcenQZGsRqosVwxXw2TgrZHxynVbFXfEn/gRrnWtYVaw6gqMz
9rIs3ssvuT/p2AfUW0NksJ9D1erujqzgXl2wz+mwXLYBmdzyzbjuufuCQN3nwGpQqEkhxZBjQnvl
7atF40Z4ApOSlcspwn9r1Vg7149gEaQ4JkJx7KT69HrEvznxJUxMrjKldIBHmdez5BQsCAxJmAyH
aJom3wLdAeHf4udwNmXdWKu0XQb8QzRYXGiTsw29d3v8vioKsQTH7l9N8hiBY9ghf5PoU5HkwoEv
CWOJyUj5UjrfpCRSpQ2lUsozulHX60rVd5UhSN33+XPlDeD+3bvzwTXyrdXGr881ofY6QKlsmi2T
EYduu7aGHArZcjNCx8qNIzzgLKfkM/E96rF5PolxZeUKtLOmeOqjaoJvNtIYvCnauUyVQZKGocjS
hjVmsI3cHLViVV75pw5rSJ1e2pdP4NieDkJAfb8pRQRe7MBt3rMMHgIEcDrgZ49cixlm7QtV9TVt
EIuNB9IPWNEK+S2wzwzUYB8D4R798ez3s67RXBLjNo7SuSKCi0jBf6yYTQmiUKt4qav6q6g7QSn6
pDaaJywSatCIAGZrors10Tg52KIdpmZTseBBG39+cDOj0XJuAerm/X6IWvgy/RIw3gBsL0ylA4ha
uHLOJumGHr2S1vvohwLg+QZLNTGmeIM2jdGGKvcfdyb8MPHgEPnLECwvJ6gytSBWoORSShye+xad
x5au+V/RgHFedf4GMe6K/LQzXNFVpH+xC6AvnRD4lDkhcjwQaBWh7ZN70QtHCgpHy4sUctuSesYx
Be+KNpSFp3qiNh6U7O5F1DepOlIJCLYLSMPELDZ7WBmfUaz9TBCyuxaGFhOokkPC2HGBVB4FjiuC
wp7K12CszrcGBvejn35gHiU239sP/stKN74Rkzsp0JcmgXFVRR55K8+gY4S9GfdxZX8URbay3UON
t654JxyHQ6/wd6LULMKL7+A5AUeW5gQML1LJjU7HGTwTsFfS2nK2aYLw2RO/Zbf2yEUBnwXMwVVD
1gbICaTsMtOm9AQgbwXwFJmcLzZ30Yy7/C6yyipRcoLCRPLyJulVkEsscHiraN+Fa0/DAQnQsZVF
H1ipbYoWmD04J38r/Nh8nbqY7vVEPxS1kBRVNTM73GGCH+zw7esKMWbqWPtMOz8z/kgP4XneogBN
4THh/XtMDoeTPpPto8A+IeCQazMfMSA1wUS7zI1y/82K1EL2rNsbLFCnhVXPesKnCrYEK8E9E47a
VpIuYPxIh71O/YvnWCBTgUHYW3MYu8S+cGehXjC2iIls3SUSXEhDUv8Ynnpb0mVVMBH4DBvLZDS4
rBIrjJaC0m00alkPl8f3uxnFFxq4PDbT3e2wbm8EZqzIbdDj80eoP37B37QCRy0MKv5wYS/vfQmD
6S5u0OA2lvMXEDdp/acKVuhbSblFT151SBJugSX4ykwingpEvfTltgwYpK4AfEJ1vTjtHu2OIazP
qWEqCnIG3TtlxT12cmOJCutjI+U3QAWCOmSZVBVDOPpnBdZDtxKkZ1E7hefPzgYNUj0xEnTIzuOR
M8fr82oxU5ojDiBot3iW5c8NYdfuLwCLSnre1k28iouyzDFK40Xcq2Tjz//K3YSwMC7kZE1MnY2F
AGhThifm8TTvR7rSHU5Z1DosWRQeUwTcCco2VNgFdszooQQSL1/Dl705hng8c9xAwsExhtkfagh3
c2Kc+kVTQD9Q4aImxtFqGGgmGmzdjxyaO2KeKvTdo7PJe1zXlbot8jcPLsLgXrI/yMoShm81E6aZ
vQUId2FsN8DXGmZrK9293jqVrUvhgpRqbNPv/HJH2K5ud8SAKoks73bGtvJTBV4gCZ/6uHCEJ/nf
bmXXZxsW6O0SvYxBJM4EDmwYpY2E33nHi+y1Uzr71eLv/ERGDx99rB4OboVk+nb7rYiPGt8LyJFz
9ZQ29QqNujOr4ZlmAHnZOX/O1f5EIdcKd8hhj7tyW2GznNKwbpaijySVX/Ar0axSKDBTZA3nQojo
awpCL0jh8gyeZ1QJDwo+BtOeaUngmgETI/A/lYcqgW8EaQCAoxN3GUPiJ6a1MDEh4dJAfotxrg6H
GCv0m+snEjJdUjmp0NgEfFA26qDuaw7OHC5MKLtd/9LyfSoBnbw5N6oSLWRJRbkisXXIfMZhWWiG
g+7WqJs+cwWeWj6Nc1mo0p9tf6j+TCd34NHszRuNUvv3MHA+mD4A17Yuxq4bK+i8rgNyWYwZx4BO
a885ZwOJuf7z9PozZZxgLzTznmU6sQuUvmqswdPFdUgfjc8TezN7OUQipSKp0676NWrADYt8vYXU
nUfwW5EA/2ljlKRFdQinzb/3gtRpKuLlFlHB9gLsHVshsfjPHC4xxshiF5j5yjeIKhkNHxY9w/bB
FgE198fU6B4j2qJrDGB0Jo/JzwTdwYZYlVc1YN+YInUjDh96tEdYgR0hjkbhaC6Wx850TXcNZ3lY
O82hTPVjTpqA0MaPrpZL7yjGuwG38C7XGqcTDU7A9YIkcBj+uNdrCCSB3Y4Eivumtr9OKff14+9U
g2rFZNDFWS6zqumH434ybEmtMTOIx0u4Xu5rtOIBRe1Ib9VY39DBNNq2XVqZ1UJy7Lo73wTzhZht
TVCm21GjRZs7QKQxHFUT0O+a1J607j68CT5KQSneum/nYoNhBTjxpvvKBEctit+C5aqXLa50f4JN
6kVuYpCkzLHNoV3kA+2T4fv44yD+aoC6dk761+yjifI37JoRKiygN7E5qCP9KkXkfES30QvTSDfL
0un5D6RWkdoWQkS05K5QCYuRzcBPIVHwEZUjvBBQOCvM03BZBGG1qbt2Efm5HLDzGmXfc61gNWnH
kyOIMfFqJN9vhn45pwLJubuC13OACJEDsAU4FwaC1jlJhDqE1K7KfDh/D5PhWeC3uPqPIdc1lmi+
GUDEM55fGmqUEgnc5eXNeFOLeKTtzy0H0+g8kiAZRsqlZ4nSDVXUuqvOu/Hy+x8Gw2CEKH3Xqd/h
XyTF1ardt6/9XReKIDLccK2QPubGIi1EHZLaeKZBt99gNZtU+sjiD57Im+IHlfvcOprEJOOBI6L7
1T9QB/9v9Q11tZphde+i87Bzp+tvFnB4MAXZU9j9nl5/huNEymDW7YVaeCMJek/5OV2K718xM2sU
DwM9CTM1WrOH9fzxTdeF86mLVCjCDSpH3K6vnbkm25j5GSsPvzvj9MT7gPQyKM9OytkYJVSpseNj
P9n+5kE8litzCvVkwtOSzacZ6F2lRIkqAnFySoHCZ3lqQeIiEHimdfWNdMpJfok1n8Ta/4ykNZAK
m1Bc0wgaFimp6Krs5AX3BbkXmCNrSMEqpVnPovWt2J15I7tBXjDlFBMGVIPhc/lDh84gwhpDU8tE
mpDSUW9ofjb+5/iD6cijvv2Cx4AcoIKTuCOafnUH4iEo3IjqViUQxKxP+wPzoDqoL5lLCInNyVyt
PAzeiVGM1Pg77zXqCXRoI9f1wI1BNtAGeJLg6mtAJX0s0BqcsiHYEu8UKOYswICNhVmEdiUoPl8o
4u17Q32E/OgKK1//1WbpnNcFq+q9iakDVDeemAwfdhee57NosHdm/e3LB72kdilm2120sxGyAeZD
th0qmlBX40JaThd5DHbY5sIkAiLuruC0OI+LbYAiJ7+4uRAEfxi7bhj9cGh1huMK0mQpsNtb9BEV
tjeqQSoxXMoYIXOlT4aGF9CwPhzt7iOp3GRJ1b3DJwHYLByfG5/QR/zbyhOyKwxc228UEcZQ5qv6
v1X2D2StK7IJGjx5rXbtgmrljkqiiBYtIXkUvGZOnv5XHbyDpXYE1BT98tjyjoKsR2xvzxYaOeSl
hig8SY7Ngzr+SloUM7FmkbmVBb2Uq9n8qH8HQ4qES/DRwhAyD/dDK5FEwL38+1nFa3zu+Am9JeqE
T5pYN4Q8Q8AMRUFesPfWKrKGCXJpMyLlf3XxJ2eEjsjZhXi2dfa0pHc9gAnyPjpTqevdQKTlqdV+
Sq1UlSQvdvKsHf29FoL673dLcC9Ww/udeT4B4c+W1ipiytA8ER92IB5yLYNdBOnVwjQTg/66fV/s
JRxO+kwXbhjRe+BYl19c7C7lbOX+JEuNw9dSC/qkUGJ4HO+dMuQ0Q+acUcE//WnOlPd7nXjAayQX
cfKyHfNKmxUoWBGOOZ0XzagTTMll79j0v/fNiqTLJZyjc5CmkV8GMFKDWA3dz3TcvVvLlzt0ztV3
jUToNGpnHazhiQMmgO67B9mGBQfyfXrK2LjyRW8e2kah89JwYTbtwjjP7P4SIaUfQm3VJMRvXFek
7nCNMr3H0meCzkSVLnb2jL11Aoz7ILHEkhkh7gzBQcdi38Sf+6myR2TxjGeIxp1YmAGxYSm+X0tC
xRX4pECjfF+iuo3j0vpBOAWhS1dP7/vubY+266XQjHPeyxQnO99RtIc7pCup6x6yv3r4o/YO8quz
Er3a2EfZmL8WErhJoytxA4VL/uYvhoM0dC1+HD7yqevoDjJpt23El8/astxlYt+r3y2vjCQYTMYG
MMs/5Th4xDbGX1SfoyjMOJESF8BbQAEp2qv4kAHdfWBmULW9nxTFlYmSdEfBxSTBd8V3piksO3x9
29JQq3caB1L3mPXY78Ane/D4uG+N4nOIVPQQXyjPKntkQyPCrggt6KQvoWyHG87LWhflNJ+6Q7cG
PDklgCfmSWSvsHqXDQpDhi5tORROlG64HCwRq3kM7DiQuuiImVLpYd7oSru8yX6WZRdu55BKeIrC
kizQw6BXMy76lsCfJY/lvTqgj+TOuQxPwie/hO0A8MCLnM7G4tsFMNQ/fYhlqy+H/VuFcRYMN4T4
aRKYl+S8w3W9FSMUVaJyjpfwpQ5iCji4M/E2D44CTLQkPZX2u9d4hIVsekXCNCaMeMqjE2abpBDt
zYdsGr3BbIFik9QnNSqvzBAzyJrES/McIzCRA36ch0VZ/em2yf21p2Po6L3vQm6QLQ6i9u/8oqLq
ivgXq0JLFUvisPhUy/96c0uYqO8z3ucoUbOGlD8zAgjRfMXOW7H2CRIeA5FZDui9uBN3I/pwxN63
sbLqmv6eTrFcikoGu2lcF0A7oefFEApTxxN5LQf9hEf6p5DDlMVdBf4LV0BS7bjMOCxl7i+mU3fn
FMcfmhgArGgc/N7fQjRK87nvdgK9Xugk10/mCBps8eNHm0Fjf34+Zc/uBpZ3ezppq9V1xybs/Dmb
2T6djMnpwiTJtr/B3VU6DJYbS7nZ4EirqW2P4hzacXixdqveYqJojrUDXIMHSds6zOyMwW9yAZ66
4rWh32u+ufXe3GDIIg7Lnh2T+BWsmg644vWJY4jBLG/4AxCF2BEOaUrMz5e5P2J5cpwZ/z3irr6M
jKQTt3d1j//Ca0vFwrC/txWzjd9TZAVjuFs/1y5mN7QSuCyfSTMXviJhCQcbWQR711eBU5TMZjJo
+UoZq5L5uZHB1yaThdrq6tR63/aBO3QOAX7/YBGg7ysyd9bxBUzGX1L89Vu7m32vwgs2qtsWGVcW
Uu0GY186thbiPpLP9E6YbF0nruer8qJJ1Yt+uJuuDcX2vRQshN2+pBZifgkizspwp7AYvsUNY5Us
maMfi2gRpslsBEN+h/bAszm589PTAsc66B6VBz2d1mQaMMrCS4L5jAWxZDKwrhS8YZee2gYut3tm
xdd3I0iNT0NC6RV9k3uUMK+JBFUEV6XFHvPDLu3RBGDPd9Me+acipWcR+HRhHzUUV01cOHaLrQDA
PpTVupQwOF2BHJlsttRYbAS9lJtCkSDCG7tG5g2jtYtlsUg9D8vfihW8wzXAT3tFo9O5xiXSyBMx
qoDbNkiy3n6Fb6kN06vl0ZDI48lrH5D9wFbaIbTvmAxsrgZRNXo5By5gyhru83ZhHLTQ8CKL9Stu
l4tii8oeZAyb63bC/HFK+S6i3wcq2CUgNntURbtBPq98qtX3/5PywTR3EoVP/mptN/3r1W6WSEjB
9kopRSiEfr9puYsEREKTm30W25y6yBWmyIZrsB/MKvwUgtXTpr8Po4JIIzlH1F1JUeWDkw28HSKw
OlcOurC0XKbkVBk/g8hMzaFqZRyBMMQCMo1/smw9X2zS5TwXfa3dCeGLRxKUMIy5sre75UeH/wiD
ytT0wIKGKrrrFsbWFPlvrBsLqvTRY/026kMqRm/uSOqv67qYWg/yTYVbacDdkeQ1qycQTKM18bSC
dBtzmhulJpUBA7AA0TKgAwxFG5S0E/QCi9IUGQNkhQ+ykJ++/Ep4cUK+Zg5Q3N0Y9JLCUnson+Po
zatggXaimOA+yngoWTh3a0My3p6QSVLPcxL2inhfO02oZFv0Ng74bntNHHQvZ3ij9WL7f+vqdBYP
GwoGMbuAPd1NNyBrQaKTJTOUd8bUt6aPnPVLo56tJnmaJ8jihtXNEH5N3Z8N6Qbe1vU7Azk6uBTY
OsH/k5R7QgyXhSW4oMB2fudgfTGGPQr91OxfgCzT1QRW+hZoJQx6SC+pyTGY4UN0CUsjwn+A7+3A
Zq8Wo6ptBOtpypOCOIoRkUisYOt/JJ2cPiCxNlNyeDMe+ud9venVGntCUCK+9acGFuzMRAVtrWko
RgcMdbx+wivmViZB/lpRjxPgytjlIYAqefjXndfKADeOFnfAw6zBAa0Wx5k3Dc7XlQGFj4jvwMq/
KIcEFUhROGiHIj5plXO1mNQgBbqR+RWFO8sB1BuRgyOvXIBrLsZj7eC1ZhJivegGAQ6sTzvnMfCc
Hf7wBEYPZr8cf27F/1E+14wZLADt+A/6aTaqAdFVWvuEN0Afk7FpthHD8YXiNv0iEeY+PMx6B3V8
aCY6SQ+DQyNg6gbuHLWRWcpRYpjoIyq3S0f4dUWokxFjzYCQnYeixtlRDJKMkn7FU82MBS4xjp6Q
FeZsie/u6Wwur8GRcP2Nu4gS+MaXHM9jjIUyN/1/6bKiM2wdr/8Iu01filM9mtAcixxcLzoobrCo
uE09vIRLhfTcAZXcDKp9i8oc5hQllUurN6WtfIlmey5PqumRkVTiBtsLI8pWvogHaIrNW/zVsJKw
QmUDJqNvcbnqvSVfphHmt/SZy4Bu8J+3In39BfUo2Z11fVRR0LEC2oCbAKcww0DBJI01PRJfnztf
qIOk76Wv12r50o2QtAGefkK9f0OBIE+mwSJzQ2H4gV0dymEtfa13Z1qA/zMSGHVT02eQvmJxtv5I
uO59BJ2pwmNbt1lbhmDFtNFYhvIeEms7sigDEPTfO4B0P5epQ2alI9xTc65ronkWmO5PwXQoGIzX
VxX62hkF2HQp9NmZPuWl6jDb0boRZ3ml/VvTn2ouiyq/hrRC9e41o+jYhg0XWHE4hHSSmUExf7ue
TBIsu/MlAZpICFl8sy/WRw7v146TcrbtlzXVF/TVZUXqmwMFBPgGA1zJtNhJHWQMAacHBRE974hN
QNjazo0dCoy7jq/r+EY8OCdoaBqEg4rebxOxbltaHfR0+K0kGjkVFfvew6A04WJ4B8+4zbVCJ1ml
VyBZ1TpN0eUiHiVB+FZFCwSc7VlrOj9M08XXdQxqoMpp+TM03Bgb96+CSeNaE9rk3AeYEcWGl/ID
AE2I+4Rf3HwoDK3Swy95puFYqyW/GZMaNNKh4LX3tNy+xMJ7cy82UBjaBQRTlVWYR9w16lLk0WlW
nZ6/iteyYzKvr/39S/vvZHqVF3rXlqd8bHcNKsctE3cx5oGWR8cCFDF8sQQu8GW0JGfBHrqccHlU
+bME2vR1hlI38Z3393sdJn7IOYOb3DxwwSYRvR7Bq3rdzx8HQIeVbar6N8LZF/j4F+qh95qzaoBL
yQ1Yju0TG8RzNFyVjxM0+38nygMrmQ741kVXR2eq964650LQhGohSaqu8kzaTDr4YdsUpbxfCygP
aiol4nYh6UBYuS7l6pu5lRJfmskXHc1P7MoiQq5KU3sCbl+/TaiNLgZdt0h/qWvAa1jEVYL3LYXZ
6q+vcisszGioBVYPhiF2SbUZo6lJhueX+7stUxI6e7rUMWWd8oLg57ge8uGjkwXQ7l15NK86qPFx
GDgDKI4hBIi64K/HfEq7N+ixXrL5vUryPE2V9uDcg+G4oPqAN8/WO91s2h9tQNxM/xhcjOhtwn5D
Nc9smQe9eC4QOtaKyXxiibn4e8G0x9pTAof+Ckxel0pHkdjsGxSNf1RUe1/ckVDelbSDpdbUSQ1j
vHTLnQP40DZgYByWrNcC8/87v0Uan+Piw081djtKHblPRTMYAaJYoyEqyiZvXHDn8wVjdYaeoGyP
c2bjdhN0me5QgtaO7xl9aKz07iqJXKIoaYmBW3/SOutQqB6vV8pJB47SqEkx3eWEFWsCDYEbYSdL
x7pQJFDcSGyQdSTZioWBM8oleeaK0CYvRYe8mTxZitY0MyZjD/LEVXgaw5zxZPXGsi8UTBvFiPsl
QoF/9lN+x1Kl0KJmhbfjr847la7vU3A6S9VXvMnr/Sxn+x/2f2aRWcdxYqokm3kYAR3eJrzdqPJ/
QufEJBdjNYOxgFOPphHf9hbk53LfZVn9plPFr36vk/2nPbEc0BgwDqB0fUmSyOSFsc+ZG7lebLlL
6U8+xn+kyTISjaXh9+RlRqDA0uWeDUshtleZDmgl2z+3Uq1pP9heCrmLg7XcCFm6PTCWAdXcucHO
HUR+woGSM/+8VwOHFVh3rAe6mlz0Zk+VvOriZXXkcINKmAuu3UwU/YhxzhWFqWt+UJdPfVRKomYf
XjJdT56rknbmWlT6EwBhNuiortSeC6M3MrKLhJZab2soutDsIDW36hevqKHysisYpDMSoBbTiNaT
mFnGZuNEFEUkXGvDyu7pCNKDOEYS/rppw9TVqgfrTDeTXTaMgK3CuE6eAMA71C83O+LHICYbx6eJ
Ae3wRWIlgDUfFoEUgIEApYMuo9EOlgD7NwmnV9o+fEfVIrtmz1D35nd0/ksxbMa4KMjAoopVM6SD
Me+UPqeAhhIPe9KKz9QAP8BLYFso8Wav9/s53BZkreewRuxzJ73xlCy3px5TINY2t/lEd8AHAVIX
FZp/HS77UuHKH95+eg/TsIkcuzcnP96d/UhbRTbw3AqiOGTc4Su84wkuRCsmrwsuYz1ftVBAMUN7
h12FqMqVfV69JmCEQivpd34FeXWLiavWuaBhkcHQ9B6pt+xwTNnnTZ5virpxxtOg2D+u+An565v6
3ZNXjSfSzV9wHVxW7m8DftPSm3+nTL+qGJVAjgcTjbjMJfLWaA2o2fK4HZ8cBBLZpmQZPrO16Iik
BcdG7HaBfrfezjSgHYaDnN8rOVhakiXXdP0Kor4mPTdr7uTKyP9siXF3nv6Keqckp4DZsMCQyqZY
ikV7yaO8iFlipmrzIlQYj130J/eiBTrnXEWzrkHcIiAeK1U5RU8KQGdrEdYooUz6C6J70e7ll7MC
cMmoXc3Hly0P6NWZ4F2PyuBDxPKTEJqIKi6dR9MSvH7dobZXXSKUI27sfSsLH67p5ZXDpxb4JuHy
jGJIpD8wIXqXe4KVmTa2YxnDnA3M5y9YMesMGvc8vRRVN+EgAF76QYmfUwU/q1dhOWGCpOf/kEDH
jhRagpSgfvmCjk2+IOFxBOPePz1kQFy5Tx9qe2y107t4M3SW0RsT+2C7NzVMlGm9+rdGrtGy3RjS
NHYZVFSuswNOMk+cXlA0XmUkmE+GHf5X2tF5h8Blpi6NzQYust5NUSr9u8f/VPFexiFCiPrPrmjc
RQseBpwQBT9y/PUvjCWLUt0v4k45MFRJ/kaCd3ZWM175QWdwqxVXDDg+XW7uT/jbblIypPswrONF
7DLNEXLCxw3wwwkGP01GNdIPzr1bVHEMR0AMhBYX5G5fbdG2QFkBinjPS3U1WdK8bAkrPtmTBDVi
yS1f7zFrRBzAvUPtHiC5/ZwWZDKE+erbQdoILLf/FXZ+PulONZkAFiferQfCs/qgGH5RSEp51OKr
Q9NsLOc3Xrm/KlmJ64zH1np8l19N5eeALNGL99apKLvmvockHhHhD5OFBkhqBCblYK4EJVKvsLyN
66MBRRmBrWYoW67HKF6UOMf43TOwS2/xYpCAX2pPoyCyAm6iEh7jXa11aoTpvcnZJvp6yr9ceq+2
i6w6y5aRotVYak9KTMvPiuEPwvi8QfyQdhyzZ7SRNEXNx8YBhqL2trmun/wSf1RT/M6RhXVain5m
xY0caGTU7WVc2xG5zA1NJpsyk2VxJEpO//RklucTCc3T0G6uWEGra9qz4l1eDQYefQ/GTKM69vfh
q8kkPZQsdAxxU+R1o4TzksYsgVdL2TH/QuvEcEI3NYcDWVXu+koL8WS6jQ+EZrpQGjPw81eWRRwt
hEHiyMbnUtVVui3UgC5qqXFyWEIkdyAZnIK+hsJXTCjryZ2XpaHsuOIp12m0+3d56waWp3jVt0MK
Mz2gC2IXwYeDoasYw3eIWkcrifPIymlzT5ZyLNArkR7gWALsiCZZ5gVZNHmBmK5TbW8EDvUen39/
aoxhUHSqiSl98L0XulMzfjtejrIqN14+5+ajXk7czs83gA80F4jKWl/psLuK4N1jwjDjT4UCy3Tw
P4zU7qSag2ma5WXsmOduJ4UOj/YWML7mVHYO63d0k1X9lbRdVfDzqonLs83zQsYha3j2cbyB9CWE
qi4QS6nzlL7gA0mqtmg0wyCA7BPIwT4sOY5sqqeVAWbmfK3NmJcwy9FN5FrwWLeGJk9pynTAFF2g
HsvbScBDYfpxqPEWEMe2WVVw7wEo57AOeNFwtEKjfQzFIM4JWSG2PvB+oGQ7RiLgogfUp37/4M0m
b1fdF0dMpOE1TVpWW04ZAteR7VxMrF5on7daQNPZAQItk+MvIQ42HHU02fV2J+5ldqaJ8TPHCFqT
y5HzAQDmfWUWPBPtJ1rUtOP0Jh+0idw+RgA8sAK6x7iwAi6DdyuyvYOV1ilMSkb7XrnkpK0uu0uk
0DvimA+2ESbgOurvu4Q/dZYSVYFQoa+Ansm7GIKw99MxrCDmGYHT50WYmA1tdNufUGxg/RB1UMkE
T1BvFx/LrVc5i5C2Qqg6bMG22AF2LB1o5+KZZf/uiPRzFK5QeTIrbWAYlzuzCdI7WbiWUaD6dDnC
/iznZ2453SyTY3Mp2p23oezCEIyNoZIjVVjZxe3rOFaIZgqxOCfKt8zWbAq2XsUZ9K77zfxYUFKp
Xrwx0WIjiJdfwjJJvo+D3J0ifJ8BueUcrTNkXaKKKNnga5XCAQzrv7BPOyYfQAIzLoYtpJHynKRu
1ecm3NHEhvT7Fs3mHyYkEbCLOGD/8oDSHwegAGbY34/P6wyW3rY5bPd94NTKn1/YsRpyZ5LYCSTY
+pCJsZsfopu9tQQYDPSEnVXQvLXW35acL2wKssx+srjZXqy+w9hsgcavudU7jsyB9SsUD7qnXUK0
MnjkiJw6hcu5HKY91flc18EHQ4CCSKWqGfcKT/YpOu163/yG/6IVx/pxPRITefYk79TAd7jj+iJ1
G2YFS29O9DNRd30taQfMbC0mkDAxoTw30M/cGwyCT96bK3jLGXmevgrvw62BkaGG3JRCmWqeSvN2
DBRGsD8rTZ5rGEnhbAQiBXE67pYBwLOZAeAnjt9FIkhbACQskW6juBWZ1mXVr5aC82AblcmUBGmF
mGeQaVZ18487KW1CIdC68bOuonTnBsgTi8YEQH/jqg9a/8ivc+eUik81s6mwg9dKsoOsF2ATK1+F
xEINh3HXSjbzPgi1NE1Jhrqdw6uRZ+BdNlSU7mW111hIiwODlknk4ulCNnqiRwlxzuwkBHCTkUCF
5hYPdpouIx5KBsuFbpymuJWuJC7T+bxIbqb2nNPxnoobMjuKWjZAo3N53YFvVgID2u5OwUI+1Jnh
N2LamDFnDGieKzy8TBu16cEoKnhQtbtrrhT56oFbID4/7AejJq4VyQp+gABCVwJ0PYall3xrieop
C8Gf659in+N3WLaqtTTXTY0gWWGSq72bLC09pnQVvdEECKwWKHn6/iIRNpc4GK+0g6xX+/cJW9dN
3B05x+2tDtCWvpuDnNUzYT3zjjAfAxCWWXYwCjHBZxhMLzULi0zQCi71Iw5su2I9Wj//LikPcfqR
/tL1ssKPQZuOTIcK19OxRbn9yM8567ysQSARSWKwLnhouiZbUs3W5GbalTgi7PIrSAt6snEsfp7E
QCZIzeD/B690KTcch/0zySB/MDIJb0RzoTLMrOJEt0gmDzILiOax+1dua2OiBAcClHLdR5MkCkhc
VjmLCz1z7B2AdmlNETJ9LL4yB4+V0z5AsbHpvxKEBLuKpTlTNm8t/fRWgPgY8jgpW9Mn2qfQfP0v
B2klY0U+DegfAHCdN/BgcC9AqlxVc9Sea3cOhXfYhQjvw2ZvzI3oCaeo9Qrem/yOPsavielxLRHu
WsZZmM3x/YITrAI5pktMVhTrc+j+yct8rDtAemDroxBLWIYRR4KO9oialVk3v5B449cIm1DdDrRq
RA5h79u+T/b3eR6cK4GzaQEyH02IFEWV6MjVN1YQotfIKnn8yIgTvXmJjO1qRgiJHdrH8CHKO0tL
FnbbZcL1vT4yhzRNm0dIj0Fg1xUisd8TJ8IvV98YO7Joq8A25gdjJlUBiXB2GDM43TOk3eqncJA4
ccD+JqWiNNmfuUTLfYr9DHN7aUM+bxinZLe5JGX78/TzKXatJ/EoU7/qRCyYQJQl/7jk0D5Kn6kc
LYeMOMGHlOcDqdpN5r7VEE0fqdskyAEfPwlFHmAXcvRzmp1fHvq/PBJEuRQOa7md7WuDonZFnzHk
Qhoj1nkcfRflGL0oZwEZ6kgoV7DU2M1jzEXZjBGblcZoK8N92q+tuLIdujYHfjRMVei5qkVNnVk+
S+EI6Tu8ImoU0z3fhjDkhtNyGqqByzM1OWIZ3NYRcvxo0UI+83DQYgA+0zMdyBVLBbkjXEEhGVPc
rUjsegCn8hWRT7lzXrI7gT3XGepbATHpKclZQAOqiROjIvkO2u0RJmMI/5ickwFEzk3SiK4l2qwP
orj1Xilhtq/cScq5f8C2ghfQN/WV2UJNSdotL6hUoWiJ4tpUKs7mnc2F/qpP5MPNeTZlzmczG8Kk
tVDlJwBUxLoidP6xEm1IWABBWkhC9EaEdSZz8uUpi/52I3lOdBCIIX73VZIs0QjSvyFeLYl37Htt
gTBwxEhC9jXPcwDjL+5zkOre4WYROzZ0uVCWoS4v4Ob9Nrie4NSIzIvKKh5wuADhGv0XLgNT+6e6
jIoFvnL/jcPsSlIJKpCpz/Pcn6dyVToeH3vmRtT1luVjPJVZ2TT6AfoRZwQRFAlAmci3r0sWSX2W
g0mGNYq1/6wBXTlLV7Xi+9Hg8RS9fOj0slzOggIYXVuvsyzolFDQvFvVaQMgQolouU2bGdVlKFiU
2rZfjRcZfTT7xwnHwIknfKQXrC8vNwJ4izRs0oei/dKPIf2qy9gPpjZltDTw9srYwYq2Aj0ZBGC5
llGJlb0bufcz4ceYnOHv7HCaiOpCaNyjEtXWZoLox9V6EtUbqK9BDH5ewErZ+1KS+g1ANKM133Z2
PnuSaKnhSVBzx73ZPkIf2/+36XfpRaRyP6V/szG1VKx6C6BNTWcU9cMlS+g78pU43kZXYSO0blIn
QFWajvGZTvwuwh1yKinmDvq5d9LXUu1wZ6VkFkFf2otgadfzPlTHluBm2JXhDw1kOI3N88VGVk1r
5jeTMC17XCQ9qJAdoNe931aRxFHbaYOUujs2j5xEkxD68CNXDLFcT0J+lYEbrjkKxpcOZEazZJgT
VZuICbcObaFmSTqUjGV8BXsnLZvRHVMwJLSYA6un/Eun8i0l4JeoPgVs8hkcp1JhUAbJP/EBaQpO
T3tjdFg4/aU9uKKqN5767AC6i86zhuZHEpLt+E5SJXTv0CeaA1joWf1/fIfbBg0QxJfkcpP6Oy9E
FQU96ZFedWhXlRhRoC9PboRDMN87AtpMrzaOXBDHYu33bH5k9EJdhnDJgHLLnkAUfvJD1fGC53Sz
4i0WDtMZOKb3Few8Cd9ElOEcwFz18TkS8Z/LonQ22WRkIXT0NTH0r9g25CTy8EnZUCwgibkb5vt4
jAu4UTRa5Uholivp41iB/1c0Squ16oOay1BxyO7H55VSGf4acV7lUyqUISeKyMo9c5FvoAG7kQ+Q
p8ApDW1OUwkIeDAhCAdSWAn5/ZcIj1D20FjnRgGowLa1MqVaGpl6XNok0KWQC9PzySPy6gHmOsDr
D2eBPVg1TPxd4jETm5w3NutJPJ/9r9QeCp/33X3kzLu7skElboAU1JvQRn/eNAgF/nCn4gKqm0Tf
PTCuU94ILkXtAEF3xHB+FXasdCBnjMea2KXlxTMROK3WHBADakIqKS9PouuT+eELweHVZeod/ryG
oAZYWETa+ECLG0M8diHfRwOCwM0N/pK5LgJAf1STnvgtfK0OKb0OmG2pSdcYUtQUdoZAtziqBF6R
BlwUGMqDaaqcIkGzlLjRbzFFTHoCCrqWl7mh9kly2NJKtu/VU9kqmzdLLcSJ8dC/nJXLkMtwh1fA
LvJsjp0qCb/Me11U4GlWLSFZSpYB/bE/WgEctrbvwt3cIZzZyXSoNNhFuzoT0RSBP3VFxDASTSrh
tbi8evPO0k0KLkc8Fqg+G2zPFqfIlmeKuxIe4oyaPvXAQVv6HUgZAi6w+F3HUXFhDK0kg/UTucFy
ncfLBvmHvcPj5+KHmiQDAUIhA3OkNH3y7Zani6ZOcE8krHby74itj/bILsQYWGv+PsATcXXg0K4R
33QN/oV3JeUVehgKYXySIvYbi7MWyjuZzPgJ9LcC0hjlkCjMYfOnMhILrDyk2MpzwMHL+8Y4kERB
kjWETV51Xk+CKXF5RlXxWFNogteUjD1LGuRo+uiYSCTWAGoN2XpppNt4Xg0XXyKj3UtMHEP1pWnQ
EJpLhsUSIh+6t69mUd4Dtekdg9kpCylonxG/YqgnQFpRnHrbyZWM/NW1lIVmnNBI6SlgeNNcfyR6
xB+l4jC8OfvX8/oQvOGutyBTp4VK5LaZkFd4jjNKiYaN7RTig9S2KhX/tcTkDcvrwJCR8wdUuTNH
YW95x5NIWWb0uAHDgaZ+wH644MFxYHpZk9aBmr1JXY02Ah+LP+q39mc9GCcnbEhYL5cTrxeGFHIe
4de0TyRxrUzj8WAVh1wuWY27tFr/7lC+YtWf15rQ7IJqrGYDilJUf8073M3V4lajGIdx2m8pUAdE
GhSLjYZdV256ueLwf3hlxlBslvqK9+bNl0ILOJ1o/kFdihEikuuxOEKg6RaBnXj4j3KV1jkM5O/M
XRFju3SYARPh2Wrwm2a3GM4lG/8kXaTf/CMhntcxMNTyWCh33I6/5GT7Gmak3NzPoCNWIfgSTK+m
3s1OEYUbHoOSqGJY0w3yIFMHe11sH/RY7rOyX2wJ79KEIawfH07SOY1QSS6OSvaK85z7eK8jfC7c
v65+VCA6jkJicniTX+Hu/D9ocCSvShvBLTpn4lcAFlj56iFeJqjAoZKionchJ/i++Faffc3mssxy
LbMCGbXOFCf8/hwhF0g1dpCw3IjBeVC3oxI4DZwhdUd9K01WpPhrEzh6DAc7DZtk4D7w77ZJZ/4X
h62i0thCiKrAeyci4Qt26YZdMYSjv7wgd/9nOWp3jjRE3QSl5cjVDsYMTunkP9F9nGYJJEO1EGHA
LLJz9cHheLuinFAU1LSMgWyxTm3FaBsd/c/LLispB0GmZvJlIl4OSOj96I2qoray/9shHLUGHAem
vHiysUJWUvFvMWNf5mRLi69V1YK7PcmhWGHQwN8JQEqEhtdcFkhxu94cubexFadCLY5NCnQJITfP
yL91bKrjZXYmhaIv60DrXOVnHjR1uVfj3KGVk/OwtllbPnvJ25NI88K+YS97oAs6TTirP80qwwnR
qpjXDqQ3U+x4nsJpncrV4U59F/q8/Kcf+goHbj1zsEomjjCdp5dOJuaptI7RwQUexodDr4edTdU4
+jw7BDE0C12QUqShh3bM62m/pfOq5Lrd3/j7lfHdEUFbD84zGpwesKRVu0wkse5jsVpTIZhqtlUk
KeAUbuMLIcja71K25ntsfCnNph+3LgciySrFlKMtg/EKCLhv4dM+bmn3L7WnJDp/lBPWTjOphtkE
qE7fNy7XRfhsPexfsPZWxWHxMy739EM6tam1AY4aCUNeOzXNzxYhSQ7aHI6C/DBQoXaVLdfF2dgx
FnlZNGFFhYTRA9H6mjjjMUMLzByhcIHOtHN/zQ6mmc8SrUIoEMGiUgEOVAQb+9qzzFn/r2YURHJ3
OxtoI0X3V3wDbtC1VKs/5O3bySwLjKMAZ2Iia0xnhFsu9zh/Fzl4WG0C7fghXKrlHkRh6SvIgKR/
Dtyoxem5wJuJlV9dYRzgZVTpOF5281ozF3MbmhAfaif51wNuYdgT7lxKgB5nIIpScCit+VfLhfMP
eXAh4hG9Viq8yydBfUJ1YXM6N5rPjz27di1zZmG3rS7/IOCUtYiTqEoDE3n0b79IE/i++wZc9yIc
bjrgHR0+0b1b2XY3uDmCIjPCvB9HnbuXLAoireCYbV7KFPUSez57l5yEKs7cGChx9VOsZAd40BoW
7m6kkwC/5HfB9mBIw7tffupZE8peIKfW6wrDTfKxcqkokXa3wZxE39oFgSUzzFm91yOb8p42odQK
FY0HkNLQfGUzBDre1Jwl1fGhkJwvZajHlUQ39FfVJ1UYDEj3DYzkn0VhBDnJhuiqLACNNMSxHAGk
D54kDTqRHe2sJ5mQZHJ7ME/U3H/RJoWQP4y1ua1UUVdytVNr2M3VzBsz2zpTRcuJbhUFzTajtQQW
G4ZPiv/t+nJELjVBnhsbqqoZuO0UySFHKve4RWwAuu7nu33j3BNzw7E0UlEa/dLIT0xo/9kkmx+4
TWEjJHPLb6D6ySk4EiaW7mJ/GwhQBHtd9MXgcb1LXPXDyfRtn1N68ghSJRbdEviufRLG7I9zYywb
ohYh+sPW5vEX8QIDlJFSAch0IpsWDlRUX81ULykvFD3k8Vlf8BRdnACRc0bWwDSpldSQcL5tmZcl
3E1XLO5mK9UC8ZDbysIu4bT4CdGllPMmVjbrsEgWgk0xRhC3x+IrZI7aK1+sJckqvPQ4yib4tE4t
p+630IhUwVAQU4Zqhw3u/t/QNaz1vrcBDMWwfMbgcgSSeGZDs2rftGv6dgx+HMdSzxImi1+b0ePS
SA0xJazmZwwZmVoYYg96wd4sAbIW3vQPqVkm5fHhBcCArsD9R3ht0RLnGlBnVG/JFU2ekhbufSlm
D2ifYKz54AyDklxm4jB07IgZkyhSR9P0/Y+wth8WYsW6Ctk6bIevnoT84kYcDZzHk5K/UL9uDkZk
o9QEnGuMTKa17gJ2lM4zVFvFL3YOsBHLEYS5irVLNEn6wPnzChlI8ras9/+FEIjXuHOsfaL8LCi4
ZeohLaD0ftDFajusc7dYOz/cwD3huhTDC/CQRxBXOGn2LxmwiNJa56OnclpVN2vWZSnRgp8yAMth
MU/heM36GN3dNFMZqNdhra2e2LW4kAR1eP+5lU11kL6Qo3/+clqrHXrpNC+IudOe4stnKYSIEuj7
Hb/ZHtaeqq/0yq/M958nLQRd1LQyB26ScjMHs18gjmXEhfi/osPRxwIxSuVEAEWEy5yOkm6Od1Xp
fifeFDfBKRw5Fn14XHZDYmNU72vsbq96ri/VIkniXgXjW/SEgFYjRCBwK3gwl9PRmIeStabf3yog
8C9YP9vCa3F/2dVNftc93Nx4shy0XtfwFuN/WW0/XDXNe8OLs+oBA32EU3+4OVVxjo1ulWc92Hy4
ISAeEme7lP1mAo/NFDEkQWx/2tJ7V6jn7Cown/S09gbtIAWCFyVsihnMiJ5kKPYA6EoRp9rHdxOA
qhb4PxUp4LdEq0XHVu8eQQyLtB7thqERVRMEMHiQKKQ1QdWLZn8oETBiOySG2tLWH2ByF55AGat/
p+yRBEdUlm4CezVrWsmNj5bjHzF03gHtMb1Feyw+Huza5xupCBQTvJ+SKWcYle6jGdR1fnUi1G0D
FrKRxBd71Vm75/FQv5w8lYjcI3Z/FgUS2RoCrJeK4QO7yMj0v7nn7MnhYNWSdJK2P4jJu6og3Nnq
Oqa0UTnfS+NJtbmGyyUkqAHdf6EE5HPtCCtStoqDzSNtaIxacI6q4yeSRf9szca88asbWY/Roeuf
hSSu0OaIYbe02x43IlK7r/cAEDYGYfetHfgFrd0kkRlYR+2pVjRXJHxhNx4PNaBXXEwSz2IPUYEv
RNNSFvXN2XSxp2BioWWSbfRv5LaRJB148wltLhdVEiEffXAxSNkDrcSz/1ijBfYmxGWapLX8qMg7
xeJ2dP56hCO8UkxyzVdCSGle9WacV5JPGeKdJNhvkMfw+o4CnqtbaH1lnxE1PDV7QjVbiXGCvIuM
BYyo5oB+pvixag/kn9HBnJNxtGqf9acCqcnjnxIaHiRX1ClxNRkrrSkawyHuR0Asd9zVrw1y/J+o
EegBG7TBCNAt0PY3ZPsUaaQolEj7rfwsgiBXk9mCUl5KRN7a7+d+zrFgPElbLMBEYKlk3/1ZSmN2
V1GQNxMKopJgrEkjGy3C/xyaYTafJRHvQpnfwaU9OGBlXT5zSHEVucJ5egpUkuhN6IFgnG/unaY7
WJ57ujAaSIzFQTrLzoAUjaHqLsds3N36V1YiHZ9/XDIOelKKsr4Brx31zNtjjpr8j2Kkd9mOIYFS
nYOtnasJ7HUp6HcFduY1TMPjZiWSLOI16AkFxhPQtCOKQWVKyfZk2/mqt1Y4yI+Dd8S3xZPPXsOk
YJzI6foS/+Bo8O11UWNyg4YKsf6+bUUKgFjUF/aQvzJYLuiXleAS50rVIK1DkxA6uV5duZlLdryH
ugQ8N9GPZJj90YI2G6CBYD6wIjzGtyrz4m9LuTOUh41sQLfgOKvaphOqBPNXAO/LDg8AdAEKpVQo
edijZiWM+hQOIss+ZRZTHcyrO4gW0sFYpTfHhWN3v3rhrPwTj1fYtXmy/zaMIvtpaqHlwhdtIcQw
z7X1MCnhhMlA0izyt4jNV6yhC5wY4J4K5WAGt5u/ZZnnhu7ZnaQhQ7U1hdPTIr4lKkifbf1qq/eh
KPRx7CwnxApkSD5xfypvY9RVlDCw1jRIVKBsNfHSipC/XBIldCRIitBIZdsjttYqDfxo8YaAy3ax
c7TmuQynUAqQBPQ9izbMki05rXrDa9E1wqzOIBEtAfjsneLgEm7Yc1xEjrXg3BOe5DyEnddutEVv
1VmtCG5y31WAeS0ZFFXF/wwdoPAvecDPTc/2BpeGLfJ9fiCgZcR7maB6elr4kz5LKVaFmQzkEeBP
Tu3PqprbXDlL3eZJZAm4B90J0LG0zezmPZYNRYBfF8pdE27yZVUL8N0f8wxS7XM0i5pn+04NJLa0
Ux2rIP+jcf9zX+OkFV6shbEgtWOahmzqphqOA6TYDV2f4+aHegbeFJkJpSQxHzMCS9uhWqgse94C
Z0zYUqqyIzcZPXpb91vwt8mqf6ndcJm0rGjU2dVWFluv73myu2Pxv9xy/0Dp0Ct5cRExfJbSvObu
dk9OqWnRpyePmR/3OMenH5bj6CeOAYF0nx3bTGl6U8MQLipEQ4Qb4UFHz1Z7bqA8wnyDzPGcSo0r
4YtVOSMldDhnV13CZpyEwaDvsxS+Tv5oxgdT9KhM2GwN30ZnHB+kqb6LUteuFvXz8JwghVWCbnfi
kckANtVnDMYiVTOu5tUP3wQgLReLTMqh4shS5sJLPsel2ndWCHpSwPn90bi8F2MRn7QC+NpppKkt
wck9z42mGYd8VfwQZrK9AT1wXsMyfx/0osEsBEAKjA+Yd7ibUl0qEtfYE9FG6aEQs4g4nHE2YW9q
3Uib/EUdmEumZEhk6REr27SXlPKnv4hA23jGoDdC987+q2R+WTo3NeD+Iw2yvOohOMtU44RLMUfX
tBNX4TH8F6hmzbIY52l/CE00f84bfgS7rUtMAgtp/afRxuPt648MkFAFB5Xz2y1XS8J74rtB6at3
uzJPsBgs9NoqO6CX/gWlygmEZsXShxQD257+F15TmXUbOEDMH6ZCkkt7sT6F4HkLITs58Ec0bc7v
OmQCBR3BIdj7AJr4ZS1MZVh59a3kVvgIfe1nCRst34qBX5PWpwiBhETXe11MSKMT1Tr9Q0Dl0lRj
da3DlJdbtL25ynYt3YO9+9QMHOSKWxrUh+NZ+molMkHpz3bD8SbR5NXFYI2TqJA7zRdNyPM8vQNC
MinFGt30NFoJNmTAeL2X1EBYi6HYfuXQYBNw9qRcU1V4pq/Eft+kxbigBOEGJRonkCLsxoBIJUie
Qf4EvnMA76xdwG9+m2c23f/NBPAXZjfxW5pz0BsFwg0rRH25W8ch+TeuP3aRVMrtdQrZqbFKsFs4
hHujWV415OQ0iTa9MkC1o//tx/LBS+wIFsZA3nNDp0HY/RJAfhPgaNXYYD/GFBixK3WHihDk1XRa
+V3ghakIgW8dYh16VcF51nmV8VFy4cCSLg2YzlTNL1DP03LKeD1XMwBOGBg0dhCJ5JnK4PVXOiDa
AtEygG0iBZJgwXOo0ChIbpqE8D4kCmmIUiLAWnEUpGemHFTUrcuKL779wlgUOIOPEGlZvJtSOiyC
pNKSr6btKN6Hwt8nL1/gGto3M7rx6eYc6LKBozxBwfrn9teKObkR2mg4csGOXPF2EHLBZQVlVtgd
F2NUiizzUMO0kzu6dUcITF1zpFxZayJJO2sMjUJAjb3tHnmLdKyqsAntau7aJLOxRH54RF0+Tyny
qcR04uverSnkjkd49NYLSb1F8Qm2WgVcndwfRACN0dX7I45EZKE2HEwN+RWII2j7QtDCGo2jE+Uq
xbkpQ0RPEDoIcftRaTMGGZYMfVZWaNJlVuQsOgVUU8uMZLC4KafadAtEemN3OOWwJUJs8ZZdxPcP
scXAivjJT4EEIyBIL32Yn8vMqnY4+wfkwl9WXhZRCczuTmQ6YLO8K4rEhayWDVuLfNrOgQq4MqlY
5Mlrz/qUDX6uIItyaBFVaPGEtJAAJVnBYmDzdygJD89I3HNank/hhSmNhe8wJDMupL9FyvtxTR8z
Pluk2hIpY0npPNyv8Nx4PcIoVgt9ZN2dkFrd0vUhIc2iI39l7mDoVx8cnm6qWYevSMopoLJ6fZOg
y1Clkl4eKsJmPbb9CQB0vOzs8NH0VEVujvuj2gTcgD5F0sTecpfIFFaGkyvP76ttkZp43PfSepGb
HO+9H07qhOBpXY2lJJpFrcuAQldxR84U2k7oAEZyzV/ireOy8ROFcbSjsF61zoQ8inHgH3NRrwsj
1078RrHK/1H0xSn/GYeJYWE/5oUqqq70AetZKr6+ef0oM1XhFxfLiP0OFlynDMBpl9gVQtyNdMRs
adMpzEQplpvfN6M3msA8D7g6sNheqDlIfx9R8tbIiBHVriNTWyGL5xtWOMnJSjk42aIO62BWqGth
sRwQeAPKUBpPVk5CiGDZ/XMuSCb32C9u8o0UmZmZ53PgPxdCdgWjWSZc7WJGivAqG9XuNa85dVl3
jC8sOuuZ1kFRoKZaEf2CBvdVmQhkUOXCLn7ic/CnADQzUNwWcfu7ofdrjVII8pP2oQzJRU/QA/i1
3f17fpRq+aB6hX7ng+jo8VnXrG9atG2VMPeWN13a5CL4UygI8WQDpYHxfi10Ig0S9H60s1yHlMQ1
dmKNwxQFsyVbhgIquA5A0Sc9vmsAHY3SpFCmdtMZ/bgrtSFZYhLpaPz2vpvnmhLEtRjhlPY6B8Q9
dSNKZRMmEE08/cF/562KvQiz0OzIvipUiV5pktv3fgFi/JqHxJICuO2G2EZf3zFGnhFEHhk1G3/B
z7HjTTacWDctBGsVa+4ZV5hHGlrRUmUePn8x+3F4Ir8XpksRmh1UbGpxepFoUvlyGk9dkj9pD/Ir
PDofHeZ+fLsHVJRQXEXlfix9xVLpRNxlbeFdbwHFAfExAmbGInQOyc5PUC5MC2WXj1HynDDVeOE1
0Yms2qTMjqmjk1gB+X1nG1xIwSyflhXpKWGedT1IwhJVlpeNYKlNZB/d02CwPeX8nYOEmq6APHGJ
n681MGtr49BO2TAGcEMA3xnm+i2whe+IUCZOqvk1Xoisg4STlFlJyFclOmIDwDTT1+gqIeE4a+ZU
dHdQatRjqlWn2S2APmBdsI9bUH+HQ2Zk6I5gE0CJYwu/40WA9RkVaD2Lza+phFxnx8IZVIkvvAJM
u+Nul8B6SWCo20hkHcER4wH+ixu1KMRHfS5vjg48H+MlhHgavdSQ2b/09TkFVFm/Q/SR0HXS+tt8
O+1vuiItH3FxXpCXo8RwRqHlpIC0ssiNyzT/7hZjvPQgtBAoIgdROodu6vnGIV+yK5u4yls1dVgZ
TZF9oeHIB9DMOUAqdSnUQULkv+B5JdXj85qhOr7RBCEP04sdEzg8HiB8ne0rmUVpvoRiw3rx32xI
IuAQkT61zZdkOxvG/KbucvMgM3lNMd0gitkr/Dhk1Jd6WvViwaJvFaWvZX6edJWfqOCO7XXW2Xxs
zRTEHDR5BT7sWSKPO5IBld8NQioNCgXD6K/eDHHodeWKJ42nEkFNepyo5O3FLrPmM/XLELSn8EY8
P32sAaXiD9p6GJxx0d1Ey5ez759vE8Gpwl/xAlrsOR4XKJjTHqnu2reGRUJBRoVmdxPZAxukHa6C
WBdd8mr+XhP1N7ev3DoeCWyTFNcmjjwtxhJ8QZc4TEyZ01nwShtf7q7fbQfVqsDSCcPMILomGBtE
hwJdh6Fv7VY0+an+0A6iuG6LL+461Fik/w7IBIOUfRmFMzYWU+xSh//ydYpJv9d7xmF89mmS+Igf
Bz7bWGg3p5QfvMWSW4wAHfxPjOcJ5QQqn7hbl7n5mlnlbSdG1m3Hd9Vn4xbe9D6EUO6fktRUeNg9
87Fusb5ZEhEwFe2VVgzhcWP31K8z6k5IhXiNIn2OPWilzldfiNmI58dUcwRegQmi9GVSKZDPalhK
egj8t8F4f+mIVHIwLUmmPA6eZwPNtyAOvsW1x3Yd5b6OzZcTPzwzg/QGwwGjsfj5sNxDLFryhBAL
kCyqUl2i6hByU1yMMmmZBhJfCZlmzGCbyDET34njVIlmau6m+d0Wgjld2We8Gx+Ngr3ap6npjIGn
m6pzbmzeGlGYBSqb5wh1GpjENHvvwxaKblAffGmQpSRjE6h9/E4w+yX3ZnMpACKyEUgHk6jLMtXU
FcrCcdolKrL+MV/wxmOd4ffgt91eH0W6HqXd/KGrVDXhwIhQR1yrgiIHfeqkDReay3XnXlkLhuRm
ghY3siKM0cLR/CqeTR5h23Z3q2BqZfOwH4fGqhmZ5okeiDyWIa31g/HAhXmrN5d6sEyyHCFDxmWo
2V717FusfSaByjW6qHBXuQm1OsLMDw13DiLWaOHFiqRodX3qJkWxKCG9J04Va8pUBNgImzvWCHDd
IyrwaTtSC94Vw74gk36Ww7c6hl3b9YydQtuBL+r547atQgJGVYBj0JkXFobdlpeqiTrmexZhKQlX
CAkXvpwaxpnd5Wex0UfOaWuWoLWxhLGqzaTDESvw+Dd39P/xHylyHJyKCbnIPT2UDYbNId2j3p+F
PJ5jRrMoUw1hzCTbMB2jceLIia4F5w8BhmstgGqsBRtyDT39bv9iK10d0o02AMeAntGPbty42HO4
r3YakTNhOjC89XTAqy2Pk8FC5pBJBt2zo4VA7cG5xsSB+IjVMM3ei9YJ9qEn6NF7/NVvZlsWOE72
TK+EX86oyck4XfktrZgETmPRBz84bMmsFauQJBwVgGyqFhcS3vBNmF2M1pS/yippgTPJuMZ2Bmpt
Abyn8zUoO5nCxbbPF+E+ik+gTEnCC8c3t2kEfSSLNN61brmsjEdm7VaXo9Dpz4lakA3i7Wbc466E
t8j7u7YLPcS0f2sqMBG6fHoa1aGu7avr28wb1FkBzxlDRxKnp2eTva0Nh5O4kerYbl3wEwHk1/LZ
DKkqHNJC0Zs7UR7BCucuve6ylm/BknYnKTMk/ztxz1B8UyV5IxzLP2Wua7wNWeWIyncpTjq8scXS
7tjmxvwVacfWyNtjuXiIi/cpsqcgvt8zitehyvVZTDBH46jDXdXIfHSaZx9z4pcHbiY0/pgUYnKr
sAwVw5tTYLkkFL6VM6O1zlzqX8Tzuya9vaHoVmjWeOebJXXw9v8rL1prnJcwxZcTaOU396u6gFwM
uVsbmZnQQj2IKPutsieW6NXlisay2PzIyRQDarZKALBTwfUpsmsRJaoQGa2wZxVgYVUFEe+EFChR
Zf+zSMNdouBYroRe7BZR3CG8bvleneNbVotO5hHehNGf9yf0IwUKT+hMkIHwTugCr5XOZ0CxPePr
AlVBFPpQXBDu50nN3XdMsOLg9DNMDaZRoxduks4NhAk3h/JK94QrUPNLuFzX6AMZf+/SaH25XB18
+7cKb+5r5QVnA8js7mCmkNnSQH234Spsn0R85BFj6K2+0trjs7jsg2uiw7Lb1eL68k1+Fcw0kmbf
zeCLKvS9uq1vVben+wM+Eu8Ou50PiJYR1JqnvQVUAmnL2HH4YcJinxLfB3wnQC8qnLUF+cPcLjJO
pup1vUSsg6VHntJ1eDXAlkzhKDZAV3H+MWz/ioktrKN7EfImjEK5HK2Y50dXCpQkzXzgTqsBYXc7
ZSlb+0FFHLa5PDz42VcJLoxYRdgi6OVNYY2fhkqt699yTNHqYEq7/dh4rRNRFgXBOARHtBR4LJxe
VlhZ3BfvC0VeBLeVzB3S+0atGYDJAWdGYSpAzkJkw2E1JitHoIsnnc1WIIU5BeS/j7EDhvRI4yRJ
HlwpDEEqO0OWfoc2FYfIh+kmVX7HJ46MghTRhzxG+ly8Scf8v6uTeHKhf7MjKnDNFEscCFsr7VEt
VXLRHuzR8Jd9zVLIV8VB1tx93uExgoCa40s5PuGA0tKTz74U5PCnrj+Xc6GCLuUmRVAsIezAjhut
1ZCLnKbaI9TyL6xwpWLmpkBu1JHMpZ7Ttn7oJu3wKmaFw4p66AphG4VK28Sxt0g0662yA9HiNYsi
1YoirwGHAKBZnZaMRJ4EFKxqOhSETM3Fgk213tB2nw12YtU5n21BHSBiSzjsGVeYvGd15S2okHZY
GV146ovu7uxUQkzNH0uL2cGNjbxMf5hOiDDAX15TV3M453bCFcKAvgbVmB3pg1mWfz6OFuoCFMpS
h/M5zVcXmFn7OhNKVQq4GJ43TU5B4cwpchIw7dvIZ0OAhbd2vkSTeTBdnbNwKC3Lo/xJtwtBe8Cs
2qN79RzODtPEcmivNazy9r2sU0N7tdt0Ndmhw4k4FfKmFOe50ZnoesRlEpm6oRtLcc3tt2avmxEr
S/I0LGISqVztqrbA5M4RKFlgz2HaEzFKZBk7SP0C8+LuAop88MjK8b2qiLXx49EVE1Xc4RdQKhaU
zrOUORIxDt1YCdVPhe74E5T8RG5nlwVcJwjGFBqXZBzk5BpGU8M5MFsi57BH2cfprCFHBjR+NJ9x
v3QqrFlkw4Es/Uq3aqiIi36Nc324xZhfjge26AN19y1nU7ul2kSnrITtK7ArGZrvWao5o1ga3bD1
PbRXvghoTh6UD0mPCDcUVz0McNBAVMaZySWUyPuWeSf47ix8tJPwiByVCM+HI9VSiJQHxiSnnmsL
9nG7F8BL+phOMEZy7njELQQwk3WAzE6xIRcRs/+Vp4/JBNPeOWpYczQ+Z+qEoT1od500AxYqLYO9
dilZsKfpufQyFCAyLAg26V9Fh6B9CILxhDy2Vs2mk8Yht9ZXFLRUHQtFNLizhMoPke9st7JBVWJ9
NsctXSH9OqA+0HzQw06z1NOjSLZOQFvuxS+ELVKSJWOPxtytcxOKkOGOFDbRTPmnSvUUoy1UR5fy
+qINVKEuImAxjchGRUR6IMs9D/fX8UUQ25W3PHKVpkQGYYeawauQ2vgsqqPmHjGQKOC6nEsSxO7f
EP0xfxHjGzmq3x2WF9+Uv9a2li7DqVMlB1zhDWC5gocvs+pjvsx1VlkMuzzvgg6CD+NZU9I2ZBwj
sBwEZFHAf8cpu/U2C7dGeMfjQSXF7i8UJOo/uMkuV1nJkvlRxHpRJFl2ZPmEuPOGiGRsPVFBq5H4
bK5LhBR3iLWmP+6gtE7pPO/EooIW8/Vr5wRcTL47HKpoB51cQEtG9ht1gdfhkMd6eHqQjNSVQuWl
KTQdehtiR8k+V833xe1Uyv45A587gwA//mgA/0+Zk4d8rweLJ1tjHwkY/uGaKKNQhNYT7pGo+7UT
ibxO8v/xuOQbotfyfftzt/LA7jINnEAR3DOUaMO/TGp1ieFHYF+LCX4VxjjUHyxvmVQhEVG3PbuX
dHGAcs2v9PotkOXahgG1OwMA0kmJoALApJo5tzXJllmNv+aV2+XkpamR3ijHNUywHDy1z8ujt23z
tE5Pf4y5T1JSxnWLcWrEjX/a/PUWwaa3Gd8hNbnOxCIxWc4AQIN2hOMwpZ4rfK9r8xg1+8TwAWpm
MgLqGNFf2btH1mwKTTEu+59ACAtnxCr+G0CQjzUZjntgoi8EWPPpgHV03kUnKth0SqSb8IdkhtM/
bRr6BUBtgNg2sYMDF2ma5G50vG70F/uCi/c8XZbQOsea/Ir8etTWV4g85ytvVB/+qTLn05pVR5ov
2gdH/Oja/tMoP6LZ76DvX7lbki9yUowU79qsQNz1JeQYr/xcefoUQKefBFKMLY13f9PBVU4docpT
jsppTiyKwU2p1VpLlTgVyxVdfx3ms06BPYUYCjwCHT8ZKTwr3ngJcoRTJE+2niY5fK6jHhdIQz3Q
7PQa/UbOLZUyyzsQEvnp9BBCi4js5Ne3ipRGIGkUoJOGdASGY5X9o6Gonj6lGpoTsOQ9giXbBOM5
YuuFLwLrFhIalYtsqEi71rV/vvfGa2mpkiYzoL3Jd4rDwS1alk3xENYnGdau280U9xchZ3LAx5/w
Me05DJNXlyIfuwJkAKfW0FsWZ2R9BCLf2CJZCFiRVklc8qCONLvTVuDw2XZuHJqu0lIIWdmzME7i
s4UolMU3QjgXqK2nSxEAK705O8kx1TkNTM8LYY1EGZaBE0FhgNFzGwN8OYjUdcQIP5IghuA1QImx
hpWt+it5Ic2CGUCInhdmdn3yfny9a/FG3CUIohz0Jzt3SB9zDGoX4j/8pkkZsKpnNkx25af8ot4k
9gDLEsVph5KNnf+EiBnUOYLISUfmtrIfGTt1Hg4FbZw0DNJoEcXUoIId0PTu7u3XebErnqEpCShI
+6fMoNuBoyT9DCg3QXJAAWeCxZzEuxjyomBiS30wbwr4/9S+Tf1Am7uBD6vKhRBXr2dPIaiw1WKl
eu5yjVH1Axqci5WALS7LO5QIOJ/OpvzGH4qU+8sk/rU+222rRUqa+BWou50HLclasettTqdZFx+A
c+xsejSSzgMpxd0+BlGIpmX+RhC9E49TIQxqRuD/dl8Xi1hX16f4ax/FPAO7Kye6D6oXARnLFYS+
y+5cZiMzlNRVAFUbFU4gPlnfxlXbh7i5xdtxRjuFY/dsa1erz4ZxcV3zRpfeu0AQ3yXVmYwQnyLN
ME4koivSTuS2SpavCR4PFpZnjOpvGBOwFMPjH3FcM97+pnlq9lY6KAZ/VZGtyIPrmsLXQhAqLJ42
5j4ydLc2zrcl+nUSCYveYQgcMz+rpp7CVTQjCJc7rOo0dMrkq8Z56sfaWR5ic8SxiKMPcnB92An0
xbj/bwyJ2s6eDdyT+94537xSewrq5G4vfeF8UrAXLfbNGz6w1bMJ8T1e7wYwmEZjcAiayPqVXA82
tD3WlF4AfZsTeZO6BTG+MUlAvHZImsImQE2xKY3sU1Im3Mp8l9vh96C13f/LBnQtZBNmmKka0RyY
FOppOj0S3AA3mBnRr7NY1MvHz71pc9f9kg750OIe1wGp9BcMNrMEvtBgQBM1MLBJ2oYVX8UqiZgy
eH9nsl2emWUed4vFrDTSCTMLlNxh7L/yaVsVcfVX+dbbcMx128hAX9uBYS3NWYxI4o9QEDb4+NPN
XAmxz6fOKdivUM0ttR0lgpmMl9M966ewg/cc7w6RKFzBLnWNKqIfrFiEE8yk+PKjwK8/0SOyeaN0
t4z4IbHDrFoDooaWDt36BgxOsGBDKevddEU1XDHLN87cMbxuOiFNM1nMM/Iug8edYmvcd1bk5fbd
W9XGL3htQveU/UvImv7Mub4cBTPe/MJ04gXzMhOZDuD1VLRj8IGA9qfAgXoOshFIWdOUTbLJxyEk
NHYjwwsSQutOSB53AWICFhnu3B1yug4BmbFSFXkA9RxW94o5RRAOYXf8gJNa4RNfZNfwRCj70b/b
zS9v/1l5rCuOz1R2Oea2xY/TJi4iGdgl4xiQRZ8Sy4m6xiakFc+SfgiK7HuDUwmb5KOSINwV5hzx
kl7flaj6RFzR8cog3tN0S0KOyAavJsMmHVEsSeBBt57znlQ4Yqr77NgE1KoapxanC1rr/HWedy85
B7cS0J560qD0gGrD62w67JzYkW4ytFxAF5GS5RorFnz6BcwfXYD56WhKKUHb3V/PewtOuXk592Rd
Xkc39a2lIc4d6hARguMlSbfTiApWPjGC4Fr6OgMTkJf0rHL5mUvhWktOdDPRps0EC+RJXa98gGLR
Q2jcWuORk+++pVJiaRy8yqkYEbpkIk1deCWoivpu8sRCmmlSABRQ4CTHd6JvUzIvuXf7KC5woEH4
LILrH0PwVjludTHJfSpEk1zkqRyBaxozh4yrK5yhZxIqihjxjK/rsYtHcHKswv0izh5EoXDOYFuQ
G7Y3brBCBo8dK3lKJnxUpB7CrGue2nHR281TVI/hxLhzyu/SARJLZgBVy3xtmg2yp2V4OMQz26L3
o7wIaFGg/DYeaE6ZsFIejT2+JMrIT90a6lCjc8MdiH/8lgQ55JN40l3KJMan7LpM4ey7of3ZXCCH
6acDXiC25EBHYCSAyUepLsaEGovBcZhB95dwx/5CrPKsrrLD9j/66eM52eB1qf6IbdhG/bhCWl/L
Fmxhf1k3ygC2iDmlvBJhybyzRQxAmhUjKrYcbYn3lWH6MbwrXtHh5BfmaLKuYALTjsWcRIofZulb
LVPVxLtB1EtunX5xPugUau4gy9K1iFHB70bmvDaFHp862AdxY/EJfkxda+ito5V8TdWxVVEj7JrD
Bj2YyNAxtl97vGnGVFDaGGF5L8688MkVlFLvDzkc/0wJs0610QmVCajSe9XhpYAqFE7iExKbjXSt
neuyxrweyz6LaSbuPDVM9ew3VHBMdorB+yCtxxerfiO9YV4LbI3M+FxfRoaJAI138FqyNK8KN8iZ
GqaXvsP1KoRlCRnlTVqXBhT9csRuXTs3MtJeWsrPkXlV2ySsummR1Hpuu7ItiNoUFcmnkRDBUq3X
qn/RQPxsfSxO30IjQfDxnoTHV1yxRDv2XfcFp1wqtg+OZU7S048t3FiCzhna1h4geGnVZ1CedWwU
5KouUkpHvY2MdG67dUt+cHdm/UsLM1naHLx3xNjOcCgLaKEvRONOF+xzpy3Aq6KdN5O7dWz9HL9B
b3Qv+jYlVJiElvcUCwxD7EG4Q/rguEvX+TOCrXwUTCjg8KKoj4X+o8DxmL5kJaewuSaEBSdFKepN
VXVbGt/Cazww6fBfH3JjJydNPTw3EQYRT1ZGgDN1DGmpX6SzbB4glkvi9Vw1495eVcRnAQiJlySk
7mj1Nu12UUDeRKz8fFg01SriL8CYszS10n9jkDG16NywRtNNtXlwaBW17Ti0vLu9FT23PKLrW5PT
yKXdWFJSRtb1kxeWJzeTzKzBoGme7YLi2Tq3IVUdRxKbYBN189NBVB6wTJEtp1txBkvCH5Fzv1gZ
lqZpkfevuj+14DQfHZvMFPDLu+DBWmkvcmfafO6E1sXkQ92GByhW0VIuIf6WAVY7ug+1Qv0a/8Ju
yUDEKBjolQKTTVXoIsfLdLevk9r35gxizOCmW0CS/Txap1bclL4bkpcXZbIqSEGYjzuSkcHxYarZ
mqYLwN1H+NKrxzcdCH9HTbXnM3Bex7hQ44bzpiGdgNm4oHapiVMuxHDgQEubopj1dTF5sz7OHeWT
2rfzDMkYKLeBUsu8ZCHZYdpUbTKchvjXTpF+h55YLUi7mAZA0yYQN2fBN5VYDvWx/1dHVOZGyqjm
NIR1R/84STp/stru2QiFbSlO7ahzDS/hdToUn041Dc4AkjsaBBE64EBqbd76QsBnDLlQSGOlVpDG
aHv6muhjGxOtWcAz7VjFULv7O+vHtlkZo2xzNbQTEgISeiIjjb+60rhATDv8iOLCt70ZZpa4oxkq
LJ2bPtIIl9Br6TflYg51A6UrzUgSn8iSHieoR9ALTaalHyYqgwUMoDEkEDCIhvSEqJJvZrpcM3Gn
WduONOKYFM2TjjDPTpbmyygScULQj68dIJO19bYml/+buB0RW/Vz5c2RhnXep6ZyAkBZ2a/z8fJY
pvDqZmqT5t4OiC2zS9lHAXGcdHghXh0NJCxup1rEtq4q1ijKjaDoqr861YHBmRf1TX6jSc+19wPC
p1jQFjIq36INcplxTW5aRcj3o3LF3UnEqzZgtB2LI0AtlFkAOuG+xDhsdPDWGqtqI9JjxUsc8ttY
VHKNjhSiXTBk/kEjD6B3GNwOcQpjVSllqHEBoq80WgBPfpSHGrx7vLKkLH7YtMG11e6qkZ8ML6IF
H/kfpLH9Xv5+fsCrpWQ6Ru0t0d9T6mtR7e7PzbTqfem6s2UrxDXVMXZTnojBxkvDR74Ci8o+ZsOX
4Cwp7puP3+e1xWIDwjq92Whp13q04T+gDzllQlzzen1BF/Vw4yu8xD0f81PVMNESGn4AnyOVM4RE
65JHA+9wQE230jqL8SQiW1BIl3GVpyMqrTvGbmD4CEL1ElGKSokiy39Mg43B+zbQg0lTngfaD9I4
egBsWIfqMf/ZUwi8slPUCPlCTYCqv4fuXxpVZQjPMEa711vUvsOCZkBmxTj7YrvqcHa+8mofc52r
ySVdWkNhRGcAA39Eaw49xMZOrCol/OxzGSJhKpSQlhB5g6Y+1T6qm9vQzXKC6ZLNZYwOYKoxZYnQ
vvNTwpwGueM7bJ7LU3M6U8WwUH9dEHcM/00RtT1cVc/3knimdfYVvqbsCPmJspDmHqllJeOxdH6A
20wHxfdZHJMZMgC0PptV0rZ80Fy3EgfNikeG0v6SIVR0Lb37YhpG4+8okzQNgkG+hYfToWPlyGUC
OEJ7CmswHGHD6vzDZ0L8tbbdNf+G7EAn0SVmWSvr5WERcA5Ov91jjeWTWCJvyt4ZrOXnHTDWDuqk
M5CvTzlSgO+5KgHMPmRAzAsCPcUjhbdD+VtaedcLETfDFzoCLNfPoG7CHew8xi3sowLZ1HuS4pSJ
xqN4oQUDKmd346aW4nsfFmwRuoTqxV20ikYcaK+iVBXbZ3vunOhaZD9ZVDAm4NnpSdsXlhZHBvXn
dNVETaG7SGiZtRM/z8etO8hSd7eTKkXlXhP+yND7MCtOqEqEQFng6LpOaF9hYgzPypB6R971TBHV
cbBJGe5uSBGGqrrGufu6OaTAOYSuw42HHgIJaJOqDhua28u+QRdf4S0OrcGkk5XapJNVLEfMH61F
oq4tqmMx1XRsbTNiZLhMAviuvqgHARmke/6cokl0N5wiz149oPqSwVj0A0l+UNYgmOZtfR9UKNpg
94OvA46tZW1+ZiNmgPIs7cwnFLSD9B+G7xGzTXlC3HGhG96C4PC/92k7LUkxK6o5x+i6O8NjvSSm
3r4b5VkEEoqO8jyVjpHIoOE/gkOD1eqm9sJfzkl20oFbopzXvQJ8+2iROS/bbfUFvGDACX5jPcLq
EkDi/moi5/qBNRIO3xfxIjVn51sS3neLq+nmQAhUvfVwamoxx14a7ikBSLISzR+IKeqJBcDeZLXy
rlC9EUyoG0C5QLGRxW3/2/sxWrifUR+bHX+Lx7cnCVCm+FeisKnKH5uPRIDLyI/Ol5Q3C6WyL56F
+4OwU5zJfyq7BtSlEgZKRVCAOHt1V7QKovgoDnwffPCYPFdDO/dMOBsdCgHAzLRR82Ea4VWdQdod
IMYmzFU9IHv1A1Uap3AfGOSXbgIiBM/S63SnfuJWgU/TqsTrV/XbSCzkQimq/f7AtaqEn1umze36
KueS3TsmkYvGR/Vz8t7lL/Hagex8WGB/6cwbBWuuUug9Dp6ta05pRpyONPQbbFRLhQ/y30Iv2KDF
5usJ2NjvmxmoXRkOtDNbdAV33yCofZG1Yhwqku3Y7Iffmfs3PU+veW4xZN4CuFQbIBEv0bswGgfw
JIw8vF5O1ZKh0DRfzXY89vtHizr8q7ch32g5EwjjDH8VCc6cTRsLpFiDw0pXQEiWS5apSMxHiCiA
lL09pEFarnFkLJZ7O9xBYIhma7J9zujqI0fdIOwVub542eyYsl1k+6uen/YnwTXo2RAZGFQDpQdr
QNThFd1LgdIZCY6BY9+IyhOwpBSV2CCIkEwVPye/JQEnJvhxntDeewJlWAQL4idqE9wMBC8DA1PD
wKO8GEHAEp+C+KlidOuh3krxFAVqlgngG0bxi1cA+I/5+ucIJ/cl0E6pnQj0aiMYwiOIdENpZJ6T
zOR1YdbdFkUHupJPOXmLj6GILXma9n7/3+X9fm/r42l3gTtd9zRdsBPsf0BxHp05OVlrZRWYbyS+
Pa8q532YSIYzpP/GcaC0/as2raQBnxprONWMKbjZwcFZuMkf9+OvWU28H//JNuQK6Zxo/DYz1zLB
tJ/GzJ//8jRRbTC8A4I66xLoHFxs50UC/xV5ClWkvW0KW1lZ9TezOvBO2HpQXm/bO9WE629bwEma
vcvvMRAihinUDwL3JXQIhU1Pmy0P+I6zitxKyqr4EX9WaQyw3hthilcJoldNLJZad5ft1V5RVFI6
AuttMiRuuen8khD3ylEW/X/Dvp90lOz5y6XalOHwtDhjhEpRVUn74++NfCW+2xf1eqocH6x3HBo7
BcXEy9XtIFSC2UgOKwAZ0RnSnJsYqkfPeFQJcOYNWNOC8lt1hF7189tr0Th7N2UT8eRnMQLSM7Ie
wtRk/McKsTdAfPQIUWywMpprSVIp2GLN2GZrAW4DVs4vgDkZV7ahlNe2RNRDZDKEk5gsVpU/8u/9
bYCKCqwWSHq1skztMxPWeyiuJ+2HUFFGr7tWJmLTSoD9OHnLdfY1oOq0+H8qLAzoXTekdj0p0/CH
SnC36U40lvCLhRDGUHi6m0FoGBadfmHmEdaewuFSRuIF4a3eAa6Ez1hChkzKK62rl7zxFJxIsSVG
yZ0UaH/DSHDbtA8bQaYswcUh5P0UKHpbPLxkZ7mIfJ+dKMHiXEuZ8xIa5gxoNTxNdW/YiQBH7/Mk
gJrfsxUkdHwzG3qPn6+lD7chBDo3igvyrS2jybkFXDHNmvI0s0sNRglUvZiT7pw23DCGb0JqpDYF
0ftBpkweFJnC+Y9COfOpo0OB61+j52pRON+Eh/3zsQDl1edBlO5xHmECKd1W5KQbNeestoL9tO4C
lXYKsvc8Qb0w9dnKRGQAelDee5WOfMjMmZKhzacfbdOd9u4tRFAh1CVb4ASmQSBsxR79zgIwUi0s
/rYK0PMcfQJEJuNoti93kLs4uNbgy8v1dj3HVtBrxBPJJ77DufMIN9rz2rwR5iVGUFOTY6AAPUSK
FkL+cKKHabzhAxKhGSfNXDaPknyjmvu3dh6P52CHBhLtitOKbnTtV37LVkyaKxjf/l6lvZS2pgGt
sIISafwP7WMSrHxexDTaL+9wyAgX3DSN7kV9FMXaj1mijvZBFyTpdZIM+wG8gLmWi3mgtv1QaKwi
Qc3W+pmVA59tt4iZNno+JNTdlh/c8UXX6PB81BHUx3ZspVbXuQwDdbynOz5VK7VFwF0TAvCWf91D
HYcWOG1Z4GZVjKKR9H+1xG9Q0CsEtFp4MG75sHcfr2/29Cro2sOajaty1XV5AQlxuPkIjMk4KNid
6iDDgWLlRK0O6PnxBo5oCY5LtH+IB2hlI9XAE3aSUqgWT5TqQZd0jrrYhCBMYO+IdglUNhML3MAK
0rbOOCPc/n9k/gjMMoHjRhoKapabJrFf9traMzLoDOIcBfYVFEJWVYw8/TDGAN3NVa/O0ANC8pu/
UKAEAEGcI8wcRtMjOpCX6mbFLk22rhiG/4zqiwO4VWlfbk5ESzwgOE1BgRokQYIRzw5ah/0Dg2Yz
L91JqOCUnxYL7ZhVndNpUyRfhq3CnuXDmTlfR15RKlYnDjs5/XQsygJkxZ+5b5qAbRIPhhbkLwWh
UJ0UsSMVHvFSsD8McRpK9B2GWue/FBwlb44obFPsbEgk25EwXu+rgnKpAXC33s34kqEL9n+CpPUc
0rmlkCl8yE51Ou5djJEkZSRu5YMZINhazo/j1g+4ARv3nPAWIrRdcMVkwxpjN47y5EogNe/nSnxH
DAyBrawsLXZOWspI9uDn+ksbSJrDPRH1fy0X1Gp0PvouOUNPV9wzhFm0BdfxsymkG+aNDRmsacZL
t4PMf0evXgEEz2duVeY7nIMFbE/RVSHHjwFcDyhllzy0e/Hq6sghBa4DmLuzLZVLuY6ga1nosYXh
5ta+tVt5RCWLH430D6l3xiU4vLohszkmOtSz4WJjHX0bR9xiRqnJQVJkNMX/7PfQGamHkgcOmbAt
yhmo/GECaaPjAv9VOFQbfqvzxdCi1XBFiyxq9saBsHxpF2CXHENb9Sps8N0tlJbWKneKK9MSO6Dt
HPX7+TZDoVmppWU6hdH+qC9UkhuMoTO2o+h8A1ytQ3n6paRYxyeKbyN7jJlKaSexTPSbfRyoyb/g
aLO7fPAxTwGba7bcPG+lEBSx2OtVEioWJItiUpPL7BnRWFXGC9I5/PywVACCvfVzIIhjM9N91v0p
iBBqS0bqy0UWdL1AqqoM5KaHyxT+We5mPKXuOoUFyKNE3Vx8QHroQMcsI93PwFjeqGmCGQmC8hwQ
YySsFChVCQG7HK97WFg32XpvbxXpq99FShnmmKncTJxinGtloL4OPsz41eREfHu5ESpXNSMDGu6L
cYs9vvu+XOztoN7nXQi62OHPfL4cYQX2GeE9nKrqHhfwTA4IshvIFaQKD9HglJCsAnV2JuOZBE9p
2c9rJ1Rxh6HJBXShxcMY23pvx673N3oGz6Va8EeD5qwhPiw9PGitzIafD5EMEiPy7waChgV5G4wN
C9wCfRXJryXarqM+k4rAKnFSzX0nyO2o/wmiPssK8w+q/odAXAd8aDzdePVkaEdcarYeEM4OvAsH
oCIPVQxbS6pJOHvUpb3cdaaazK9LptinBKPelldTXIWmt/Qz5NuxLLUptc8khOYUZeP9V90sLYuh
k0pdUMEOQM1WBz/mhXHAesqpa/mhrnlmKtcmQFfEg0yQyj3eA5/iIbhkUy1KK39Zc7XjgAzG7r3Z
IKu3VDQmOOdUYtRKgXm4VHqPzOXrue/hClQgfBe1uRPfn6oRR03JcI428vudsvrL2+KOwGNhJo2R
GHqSfCojMzB4+1IKmC7/T8zh3VZNojQeRTIwVdQ/oEmX7Gv/kLkYA04J6dI+IcGtRcALtJZmjecL
1xqH4fa2cMawN5afuL3aT/8te27vi8Q+bp1TBW69nOG4Kzi3JSNwu0fmOm4vCJafv5PSL0a+Uyi0
19NwH5DmKo6WjhW43E5tdeh6bclVM8RNsXEtVw2Ek6XEH9QqD+USqle5Fh2GG8nKPtqM2qAwiqud
rr8nbmmKnnua/VvPt1DKpZfZDloI0DKMZ/n8lelysCSJuy72UpAZQFVnA3k+GzG5tnIPqJknnq2M
hj0cUQ5+oTPKuhYbxMvqxYtig4Wcr/G18RTFaSOTvv9r1VQOxWckx6kmOJo00oJYW0UO63AgnASi
BCutBie/NupcAhue7Pw2gQIaIP9oQU+ps1rigaz0dufYkmLtSFOr7+JeaRkKx/t7qBTJPTSgt97B
AMLdUu5lgydmwADYwBnP7lObh/+ERskZPlEX7g1ZCMdTrzSvpjvD4W8P8p+SPQBCmesCB8mQVQdx
8qGV14SMWN9fgFuPsPUiYZL8pYzqTJWiFD90Aqpc8hZ0Vmsk2UcUjPMKXJuAf7+l8bvmf2vkSLxj
XFx/VCnE6Y5reJOkxK1GPOp/zxSxMOqOsct3ls0K6Opq09b2Q94bftrMoH+EbUwkt133n/8CSGI3
sL1JXakQq/tyd1xQdWnju1Y3AjIwE+wmbO5x8i7+OiA1jidSEWMdTpnDYkyXrcmozw3QCcNPRkwl
ABlDrzK+3jNxBA8Ry7NizqD5ZewxVFqUxgMPWW0mLwvOZePfCPnFO7W3fdn+gwGZY5/oqEhlSrFh
jJJZumIBAf+GXLW3N8A3PBu5U3CajQLlgoPOjuBGPyXhgEPEikwq2JT6tyX6PFXpp6dxrac1N7jj
GGslIpQ/uoKzS+VrBK6UPTD+ZkSqO1l0oUXx+uN2sejQFNeRXu1BWw1bJkYwiYbmh4H6bBy2x4Dl
RlZnoE9uJxCavchMDAuipKEwNWIIx5EJ1DzkmjdJ5IXs1IRpqX5hugkQwxy1p90dAyrRnuYiPo7E
5rBeQ+zL6PBjw3AewZjmiSkGbWVNN1x/0uh+Nr/hmu65pzcewTHFVocNy1jZ2NjSbTmd1gt+bvHb
RuSMfKE3lA2P5RJeEqzejcJTfDEiUnyv7OA+AJT2KtZ4C+u5padpwEJh8i9nt380ibqwM8QGsSm5
CSG9A/sHb1Q46r9tksfJYnPGh90E/e6ZFAj52GuEtDobUyV7gz7XsFmFzzSSq8RelUN1PzpeJ186
0fHS34tmmCVCUrrCYUJsBayNVhII9yU5MLCwzA41WQEoru4oYxpms9grXMA4bAYt+BVBQHHn6Ac5
tK0zm7P8/m1EGNPXM5735Ektr7Z02Sb90SER+xQdzAq8s2kcvIcWkuiO/iCLVmx0LAaXjlCN/yxw
cAIieeUZQTfokxDVSGHKTnnHPkIxOa0yU2ePY4IfLatk+eVMeHK79JeR/XECjpKHFBZ8WnZRIUxi
hq1CvcWNYrVyDbFr6OAhaaIZUsNKZ5/qVmRZkTTVBQY05w6dfgdApoAtWnIxh7y5+Wq+cpuYb2dY
v5WAQ0SsrPbKKKzuR8SX0yPRVb1811FnULAGG6ghF/QjN2zBzckSO/raKmPnVb3ijUox3tN01658
29TE0nkrhx7X36QYzTP7Ugz5hvC/w0FW8jXKq4knxYpH3COEivfaZnTcUF92A/ZBlXMJXTCPcSYQ
nir2Ffc9oR93zltZC45zHqFF3xEYWtvyIEKf/BHFxC83CKIz8BnNoYe0aX5vpvHRuih7fDDBnrnR
mEHC5L2EWxPr2nznlNU/HRT1iQT+RR+YVX1VuBcusOnZ/sVQ0Tl6u6Q7FMkZgf3K+5vNuaBKDmwT
xk2I1ipbE0R6XPHWlIcpfCovipmFLQ91gBU6okuNxoFr0PqZttWKwAtv4nJ4+IDs4D+htT4HJSya
LzNu4MrHfSXtZGBjXMtL1LBVqvgVtCJUxtbsrFC1QyOxWnWNn6I23oMLmRD3haZVuVnf/X6GUhUR
iIwN+TDNJrSmpZOjiqoxQfPzbhN1V+xsbxsk+MialnwFolua2406I8WJAqtbBxHjrYDB0j+t9Pq0
b56WIojiZ7ULGcOVDIQQxqPhMSM6ki1RlZIFTTADWdQ98uj/uxsakDt7HAtKab515v5fttpzIBar
5Ka6zwyAf8oezXyKwHgpVB/oiicQrs3+UaNdCtVbheeUSzKE1UdH0deNvzWioyWISPR2HSgAiMfS
YcoXbTwW5MIy+NZuLRNRo5gCZC4IYxfZU/DoPppm+g5PMmMkdNHFgINh8ucdGJA0RawhMpIGEb7i
zuSKQp/0BjmhCzxc9WV66D/NMpT+BxFGtZBmNjxRXEfOv8Qt2L8hWkVHvrbDIluV8b7IHZu0fxCw
kEvdwvMgorESSfmzBY8NjwivG/rNr+Fb0VZdWD6K3AxqbpqmYQP8rTG30Ajm28LOC+Zq73gMZ9bz
AQzi2wIemoyCMlrDTFu2r9yseH7GEn9YWcr40lRGPh6s3s6CaYOyHnOZzkvw4LpTM7TLUEMEbpo0
T8bMvdoZjLM+KfQ0HAAiqkVN3E0mJCGHB7kGeXkx2aawR5mNRmHK0+JZrzogrmgLBhqjAN9tVGTQ
gtKOgR1VdPiwEVsVttBFOclcf2br5dG6/GOR6GPlQ7/o5r5BhFasYq7rj+5mFtDgb3VN+FGgv6lT
jQsx/ARWrt1zS7XArPWVqs9r0RFOf/lU4vdCFphTd2zY1gYsvB3WD3wgYzCfGNDGb7ZbHrOK6ReJ
lAo2JaTEatSBsly9G31xSuiTULSxCw1w3D+4mctlmKGH/F1pcfriRadoF9IiwYezYxlqCXZYSS0x
qlXYa/xLfVeur2GDsWKVzHSfV5M28Jp65KupsQLDiNSHVaLqzzLlgb81t+AjFoqrK3TKUgVqSzzm
qtQcBKqau9kiARW5nvbNKouYvmb++lBK78b+5jC1tLgJ/4dwVl3ri9g7droVsXJ7KFXcZ11I/9cA
mB+A+kpT2dj8NvQguFD/mdKqyTOz6aSYpfClnnbxe915Ox1PDkp6Zg2Uy6Xqgn7T2McZMFtEg3+R
AWoBIviyG4Ymo3RjVAmCwxXKLh0eZrdRxI/QWRycgNPVADohJSkHiXrSiyJa4yKZs+69aGWfniDq
dnCpdNIbW1WIpqk91XmwIjkCBsTmbKvvE0oFLrW989uGpsGAD4WOaQUdmmdvgbgUnMqa6/kHFwiZ
R9xnaOw/8nz8NKDh/plJVzqotyIWUydkT9MKYE9xDRt0PDe0EZlDfnXcl9YfOfSJ3wgt49FPgoTo
yQn4UZY8vT1NahTWF5nNAKQYfkocFR4Fv3KLYrZEVnz2S3/W0plbsk0VctwxHxshcv3NMWEYusyq
vzmeNdHbsc5ur+o+nuzF+uqplznLg5UqFYSI+w4oz0KiNM/smx9njJ4I9NG56edRpEZ7jI+h/27Q
tNBmEHkrSq3OpHTZEv6DhO0sNSfNMiCrwDhFyuiRKTKrDzCYwBBAhhVXrnYxtKMshtQRHuQFHtxi
Vn1AEkxreMuOF4w4b/p4pKQg9tZQ1yKyTOHy8/X7NeI69lMueTmMsp6aaVwGvXVAd1ulHYzdyTMG
y1RImZbx8GoAH1DMOjjNxXwDp70VxJT++obuvYgkJZ0xvRNjGp/FYhq1dUqPbaLwGtOSC3hjgGlz
hKQG8WiiuSBHdf4R3shzJSaYtOXGuU8oMTlXJ9xX6qlk8EkRGKf5HX5ejSIGmUXM8DlCibAOBMUO
idKl+p6Q9/0E6BivXbOFsjcXZKn03rZcoaaZspdtNr8sH3WpGRxuiBnVWmqGM1nVvFcxxfuCxpDO
77v2BVUHIWZGn72BvI2ZmrW0qCuRMPvopplN4L2lxmuhqCrNS3RC6A5Tl7B/rDsnrUMyNUXyRIGX
d/NJl0lctOAZo9+EP45lYmt1GTcAdhc2Q22Y1g+kF9RkTywN48NyK6M9V5MxuCABDiGmy4EQuz89
pley9A5AgLUoR94t8Nik9ER1cTDZIK0Yii4dzxmg0JZKHu33D/9iHj8rAwNJPC5V/zKo3J1z9KpG
t/er+WjfsMIR2EKn5X6vQagpM1slmQBl8hQGO52/xEIWM3ZfPXmmt4TopJaB6wfWRWoVG00Q2ztf
xdY1EgjiL5SUrgeT7WrYuqhZjDSFCwLqLbYmRzQ2GuKbm8vO9e5mMaGeD65qmCjEbTquN6pOGIFS
blg7tlJWMwvzkzvjaOhZzA/NiILJNJKW0XNy3MV3PSJNIJTtZ3lVjwA6sbAULgUguv/lZtNYr8TO
0Ry/1IhQWDrciSYPaQPXs+6+5NP9BToz3XnY4oXUKYVLks3GmxtG1DezJgTv2BLgDoAcFGaxtCcI
fPIsSy9Xi7NDfnOBwv3uDXwEq9j1Fv01yA4Dyz3d8nSFl+eZPGWaCSHDmTkw0sX4bAyqlm+Du2Z4
Y/iVgBzaF4aTdWD8liNfrUDYLb1p3awYwhubCMDRPPS1Je/eo18vAl3ZxEH1bmNhF+7lqvU8YbvV
3A58kjASmCI8+djztL8DWs1NDqSbnUsiFBrLXnFfpBq8XibuhylTwwdNuFzW7XieGV8hieiSwGTA
GtYc5M/0bofsn6wKjvgDWp1yvEHzHoGbHgQuLvPIv2GtHAyZOdlMxkugLz3BQyiLnn1qF1D3QKNR
XOV32gXseaRkm7W17mZliDnWViGjrRxiiDsiKRGFoHJwd43vgtJTvYrJJNzgrCohw4Dp3tBc/kRt
4EynzU8pTc4GellUD8eJOg45Q/B7cRNhloPzAyNwiEGLGX5moAgSi68lw0AVbu9GfSkUB8Fo2y+K
/3WDgJM1NUJZMDUazN8dW4pf1PH692Q996u/C+BE9U8ifF/4kTWqrKlAmX1zKJ5IgoCty+qxjEG+
Vn4sYaDnZlzG/sEaDyfPrrLidp4xYCJFbs5xe7/eNn41jlXMMewDNwE/eDq1zjQ+QCEXYDsPpc35
vpF+mGiT+bSnvd+/6YNcJ+vuQmru7mJqVUsmOyKoshtP4WcAmmeMJJOxAOMgUNYXcN+W1didnx/b
UI5evX2zNBgAWz5dQUdFTcUvWxp8c8QWqregWQbgXQwK6yIUb1+p07fyAE0Cj9j+xDlCgnUwyvOm
4MJguqD1MQUIeCTKhtgJIdu4eD5ZSwr+af9Cmnlt05lwyGgYJkmkSlZNW7BYTgBpzFA7oWFoOS28
elCC0PjQOCZA5soHQLuvwHEaR0cfMjtDcJt0TJhxZK6/UsQMbhyVBZGbGA9Qv+TXX0Rdd7XvtpwY
acBFH/jH7BjVzJaV7MuRr+jpma888dskthBhM/ZVkb0y8g9LFg1rIQyoHwIugf0bOSQhisAeYQhT
n4b2e7TJ9gnaoXJrO+OfgTpX/lstHRa8OlmjM/c7ogUEoAnlyTvj8SrJDLPJmgG1gbjrbhlLtXZM
qUQnGccdfQny3K0TMinUy0CPpcSemElWtSW02DGsv3uq/3kwV5Xl6/N5dcDL0wPvKuhrXrr4QWZ5
4KTk8JZLxknF/wpgNm8uruXtyFxD4qs+eQlVxA7GP/BtqUJH0e+otwT1VpgEXxUjdb+KFYeAA5Og
E4ghGgyupxkqMUPpIvPERNfd0/8EJnkFcLxM3EG3bH4WMBXJCdDyq6WcvjoX2XXG+3gpPpn5TWqw
WJnZy4dhidmvmeENsIzjUa5f5z09vBwu8NuYWUfdMSbyiGNBoCleOGwR8GZ+8IA/VyjVWt/+Kbju
pCe5VYEnHCWkYtPD2SOSAz8KlNbEn3v4fkw2McTOOawfVtUdkfo+GbIH8TblkulVjjosnRQ7aanC
9Ri/91llTe0Wr/W6lu9bLUXZhj/xqYb/Rzq9cCZ0f94QmxJ+FovvJUvfB60wM223wZanEiycTIg4
JqQGxuFD06sbTgINlghYaD0ecmr8dgdoyUiIZo+Po1d2Y5DrHZFqlATUo/DFNwoQ4BeCUYjSv7ct
S1bcinGvIcrQr7sHTbi2LnMHPJcJH/JcVbXRx23kv+wryJQ74mE9NpH8v6PJXC4BV7Mz3W2WIfb4
NuIIDZKcs9WoolG0W/oe7bXorZgRXnC+A36vUPQfu8jpZblGkYpsRiK4Q0BNRk5NLQC2vt0Cn0r8
bKOPykmqjxNKehBZK/EH2E3LjZUH8CstHvnhMTtg3sceHtTU8USF05/zsC54VuVUUOzHEcKrtvsM
0+vUhBWPkADjDfQl4ECjzaHPZS7bdJbV+VqqRtI0k9LkAF3N9uxVFR7g47BvgkEsHdnzphbG+HeB
+fYeSUjIl/ajygmxVQZ6tDanPPvnLsF+vEDO27wXegpTNkn9F68lyy/R1NpPxA5sPiyXkBwgtLkh
0ud3tpRqOf22uziHy6ktGQPl0cKvhJBR49AnbRjJI54FiHNbCrMA5ISTr88KVUa1IEvmPqcQ0Hdj
GkEi22bmlYgDUR6ukk5Pe57dHBq+fK2rg7WFSJUbX4sJTCHOsy46WyfYHKpMH14r0/Q9PeL19ewC
C4aapYIKTxPe0owdP6vamHEsbH6AGdHHbHFdYPV9WAMcaYeaq4ZPQWmkNw1c7p4FVp8rRbUpNqEP
3zXUcoDijDyR03fpRHNEB78EpHdXAfyDOXugJc/wvR1XzNIibxPVVWrfbAmZrG2XqmolQCh8hEDv
DJk/PpmdYu5mfY7eJuNlWHOaPaJRq4DlAPNv4IoabBIUPlnpL4lMZoD3V8at1R34TMWWHUix+52V
r7SZD8a9CHo8hDh+bzVTuZKoJ9WIdpSTVRezlkJTazyPBzdTRodTPBvQCMDN05Ni5OGkLBLoG8oh
ZxC65I/1J+q0QkssySFT6eY+BH1jvOqm3dOevJWvGydA/IDyl5vJqNrEEDctfT0FjzjcQgoKgwUE
gZYEh40IIwvj+83FPYytVT3LzTmz7qwBfJKL1XLRRYJL+pspALywhOVCKKy1MxrvbzMb8ZvxQ87Y
xqz/FESn0uqMbkNoqmOXEZgu29GXMSOmLEPhpFQicnQHoQFl8WhYZl14MCGyvWV08SUby+qG7Ejb
Gfsm3AfA3MmU+Y4Z322czFz3WAg+jF3dSk9JIejm6lYHNI6o67Drue5HHCTEvilKAhrGt1X/vxsz
i317i3rEgxoUSwXXeJUxUBU4S4lX/u9mSukfw1+4bvJtzz+jca70ZH1j8YiPZqzlbaqUcoZY8Pf+
lYxM2Hk1pphsVd7ZsQ7de6oy7h8i0ZO9jmdWlIcPprTcQEL5hg+/3Ix6aBwqMo0gF2aLlTHm4Vh3
hnkNq9voWocQYt0eJmJ+RDOmmAuxe96x1H8qodZj7MJ1eVqPYIWCRrwcEJ3Tp7Zvot+g2kH7EmwO
OT8hd3Dc0igKCWApJVNaYVuKhc+DXaHAmO2dtL7gZcjRaSIe1cGznG4E58hmITRMLC6F30SSv/5o
kicQ+8DN/OyFVo5iYUuZKJWLKmvoQuLGhpUxeu6MBzoM40BE6cQDFlxMabRhI8gVeUubj2xh/PWa
xUO2hXleKV6enODBGukdt55qKbl6zN//8HD5DLtLaVcx77/BZR+3obli0FPczTsjbXNKmyq4IW4C
BCabfMy1Znf3EbkBGHTOBl3Fs0e5lMorAvIjblzgxqXCjmRTZaygpEpD0Grhf2XBVMmAmDmrylrs
ehgcaYBHk73kGjlw+6gnIV/i88f5mPJ2XlCLstRhJF5jYBe6gbUaAEP2hBtidD+X3d51MxrdJBBW
NTmUwXs56zcWv9JhIUfDbHjxdAVHCFx7gGANWl9KebzOqsKDSjGKneirk7BZttCPqRh4COcFptLu
NwoKjnxfrVJpxdTfG1PsVjay2bq9mP6wrpXQv66xyTvS+aMhYxAAFmMq+EsQRJ6G9vbF92DZsYzw
f9LHAqv14o3AXZuCquEFk1hoZGBZso+gA/HggtTgMk4TIQFLU0RWdmAQdNQershGRenftaKBSuDv
+35PmN3RDGqDVRF8ohRnUsOU4m6sVGQaAv3pyHVj0ojqWvmosL05sPtn9vYWTEf8WbUuwWlfjGN8
oqOaAS3U1VMrHoMxePcHt0o/9BcC1QOTzOhdcO3jA0zpFy+6zOAcB3bL4KUH+mX3ZvTnIUkG4iv8
OVH+2QObh8Ntae187vUxFRfm7brnltYC+dRJ37cYqKqvtwJbTJCtdY+dkB4DjoGrOebXs3R2MYTO
IBDleNnHGyFdE9U52BpXgtMHeK8WvF/QawOsHo4YYhQ6c3dIwe0eErP6kpzllggdJKpbcDBN09bb
Imd/JpNeTd4oF5jAFgTjDopT7kQKO0QQfNIAiIExO38NwwNq73oylgTOqq8i05Gj7q4nwX+Tbof0
pYXw0n3H/e3KFh9zXJGdPVzePUjewDFJPIiJl5XeLwFnGjH459YS39hjSrPByLVRGAMy2FT06xBJ
dT67VsS2XkhgMSf6aLy4cbbbC8uRyVFvFCQCKMhDyfLAc9n6uA4VMTy5Af8vC5Ap3rEtC18QVSsa
x5JoYcmpV/5r+/KtYuGNNkqfNLpY65rM3fJkLnpaylNG4QUMxQUfGRIklHIzyGppo7eUoi1b0x0i
GgOrW2UnoLjp6ZzKaC2b/Vy51waO+aYvA0WZsD1Xz7RgCct+i+PJ13+PN6I1VeJ9MoQDaMF/jZwk
X5M8BGJ52PgPeDcv7C6IZanPeCmKw5XiqnCk1lNBJWFY8aJzuNErNoq6gGKN4cf7QpKL9YFsIh5W
1ShbjKZuS0zxydcwxDkNIUZsm0RCSmHFpkwcRyhXYRXEbeo5iDQ9GqB2rwe3+lrPNicUtkC12BFM
+BxSI756DeL6unOzGn6MyHaIecE5WC4uTKNjIYNIji545GbyUORQC20sgHN2xHR/twAc7bUHdffc
qYkAC5XWa6sEiySMnFnu3y6l+HidDZ4AyAOMELuAHM3XT/Cv0fzwvT6X8XtL4LPglAp0bUNeCwM2
OggEO/YVhm7+9puBc7VCuM2X/TX6g9RwFFXXzHYmA2qEJdeuymN6lLQ1bhM9y5G/pnip4MzHLn2m
jtoXKUqh/04A9evnmXZplQlSi47kokkf3filg9vn8wI28+brDhp4MyGVNk05LylnoQPwFnlVEBrn
sChQmy/Q0hqasZEMGZPkDmu7Z9VfkMvQf04WV2Mj+S0+Ab3CKJ96WpZPV0hQwkx8rp2Q04r+r1y8
am5qDJFs2VxBZE7XV5+SAxc3fVPo/xHToFHCmqXVjHlKKoG7NDhWkBJ/NP31SpAjhspUhQzTn7jm
K47nSh4bZZjQ2iWj2xsxQVmev22sWoNiHbpFZwdTBOi7aknq935Mjsc9YOcb13gxLZHJ2/Z/gfwk
cZCW8plAaFCO8BirXL4XyNsvmhpR+9aFRRjvYvX+znd3sGlR+0bM1CsbWH6Z+Rx4fvPcZnuxu4q1
pMapGcfzY9MEvr+VxW7A2YR4mj1JGkFX1cARp4/PbffWk2MjHlfqIsnHtgYs7iDBxgsNwhVhsVmr
0nKYPOmYV8L00oGS0jWM78mVvQ+8Fw81gp/O1QVn7SnBaXottDoZG+sqMp471kLfmaYE9zmGpnFR
s4io4/e95IeXxN5BWRg8iE2KdZkL096pAPQPNpx/UMgvreWWASxBPDs6AtRzdDiSJfmfeDJQYqZU
fG7HJUFefMOtZgJpa5iAEIDzP+R8ukX9dVAhPqyjrNjl19vmh5pgvwelMb2HCU3RpCfNPVG6eE5H
maiXmoE8q5jVnVbfg/zziFnODlpkxTo/+uL6Sx6PHRhZvFHABUQzOoen+F5JT3Y2e0Vz2IpHcgGd
jARA0zcTgOL0DLOgQrfiCb0NX1J3Vvnp++n7ymasao1lHh4bc4QOdXFQjCNm/WQYj+G/sVzOY84C
56ZPphyWE+ZxZ5HLzlcjruQx3hP8u+egbvIIKF5iNp2/FQJAuKh3VdVoNZXsH2XWuyPp7ilhfcG2
2M1qcdwExOt7IARKI2xzfev3M45Y0eLrdX3FZWv3rBopFuLud87Zwy4oDE3SjRbJlkNf+tVEg7LF
3mJZtArd9+qWJ2LSAY3ri6wZ2yowxJ3ABYGj4ccBSag98DjeDsNdwGiZR+KnC6SRKTlQ7zMgkgj7
N95PuNjzEpJRaUhNTDauFtyD7/nFQtkpPRl40foQRb6YqMk2FHCZxk3K6lcAqKNOZwJojsfmQmOi
veuplNliNA8jDo9jNCGppdr/ncm4z5obwh2ZrjL/jlrINk0pFA14hDKLn743E6WyLhxnd31TdrKm
1OGxll2ZO9bsCWEkZXchFmVQwVga5x4cSY+rl0n80YXJJnHAqF2Jw1inYDZoC5S4zlb5au6Qvijz
w+eBj5MKKCwgkRP76w/oOSizvITR5c3RjbTQgR/PklbGDFtL0AN1dKfJ0cjDrjY0E/TJ/LhQakdt
gB3epFOklXO6O3esJrv33m6375QHka36gkobS2r26xW3xU++iPa/wbBL6Ss2dmjQpg4XqUakGvZ1
WrTAa3wRM0ObrfjsrfbbUBdll8esn9Fe6fTRMj8LynTJI4UCRUIRs3LYwGAijHWndHnLn64jG8TJ
f7hJKhV/pZAJ7Wb5MZR5hT4CnTQxRuTFPzR2SBxC0nKprSNntdF+dAK/FMIXY49LIGFYW/qx/y3o
vYpZEUVgergWO0t7yF+75+gJvy0CPWLv7agDKdDq21ZpspRvyIreNpzbsFF0tjql21NBkXAg/fTy
4NSIKfvtCF5pT/XB+cMn/WtVUErzU0BCU7VcTSkRgVU3cytQeBvccK95BZ3DdIkboLozomqXmpz9
XBkuVz26AQzbfKgiMRJWA0Y8ON10BPIYC8JDL5EGHt67m7h7HQvKaMQjONT1VPEiFK5hfMFe/fg2
ieaZj6u7tmM1rTWgNvVNSNC/J0VSYebavILHDv9yIUMT3eWHkjtptK3cF9z4r4VpxR4mQPcs8PXD
wy3cQao5ayrirBd1xBScAEQhiR2HKgTcYwTTQjBYUMOuH7U8B9E/y2v/A70WJHMt6f066BlO8lJ/
SVBiK8M2byzt+lkdyPdByLx1Aur2g0nLRsOPilwlgquDbr+CaJtZQLnMFOlXqFwEudeUa13adacs
6fczoEIfds77N0CBhScggnU+SvolqUdzWUqMZ6J82uxtY3i5UkwPTwuJ0qfFWsJPbOejq8hUCTsm
0424H/HQShVibVesYB6VLp6T0pNTMXqFXPBk/F/aApWq/KWltnkRNaeLYSAQwOLbVLC4rEoBa66l
2cQ3VesXeIwBOxWKy8sLrCrQuQxc2OShm3pEuFCoIaPOv4xZQNZQbtlKRVwoEERFQV40s+U+Pg9/
bE07WeuklZtkWdSCLcptPlQi2JOHsAf0KaNqj6ys8QGiJiSe9/02mkcRuTYI2LtNVXujlQGFYz0w
caYPVmRoo4IZpx+xK2qCBR64MxnTCyY/HSSZTtZnyQVrBai0EkOnugExeyKps5TpG176ST/hKU3O
3dj+TKKrlMt689srg5ZLe5SIUMjkuS5RxnILJzX8ns/0HvPUFzgvUVVBzynEPmlqWt7fr7GG02kj
jfIxV8JlVtu+1lUbYK/IJQZovETzKvwZfRhkLjSsz23eodHGl4UuuLugc2NsjENOdlmfB8UBF0iD
bvOnAPFAL4Ya9f/amQErYiss5jwu7QiqNaaUMfBD4G1/z5l0tg9su39ydpicxeSUcvrp+kZOm+I1
mV1WQl75SvYTsLQ4AQ3zOQgDUnvdcGPls7SwYPI2NDa3P9n0DHUa+X+0gaY98p12X9zFLWbwrN2A
HIPO13MN8EA69s92eAAOoDPLOinMTJS297g5NCdy2wHovvetF+0nwk182GZ+KUx9l5oc0oSztv02
PotmCZBi1RAH9Tv2LgwFBvXRg6YwOhjevD84bueazOFfRL+YkEP+1TpDdnd0Jq7+BAzG4/dxU2+L
ZiZycd9zpl1oC1cEMxTNJSyxG4mKFjH2wftEkTW5AhWtljR7GZSAmjZk8EF3WyHN+IlAeGpBR5Dc
iMHdVIRN+5QSn/htOVeIXlOTsdpUlAlYz4SNkJaNFEXm8UujAinAGqApJ4IqzcqgasoGVF3A7u1K
MahuXl/KKf02Sp9PlMq5il94Mb7fbqeLaHrYVB1Bc8uTV6obAmFeDWkoYzpXp4/v4aoAUPZ1LDvL
OiJbVzV3BwzLjSAIYClZWsAybwjHr0jeXHCFZ1FHIpgiWChcOMo6/9IUhyJ5j0uPWH7jYgixPjNP
1K79vOwxZYfXyj04/MVwwgqa0VSqqBRBK+RUqK3YzDK1WOgcuovIGOZodDefbymFz+GHtaYoHf2G
WxzejG9KiQEjCxNabSW5BXlDLUajTKQ7bchqMsOe7Ez+n6Wo21ktDP3y8BSja47wWgvfTp5HBSIG
edXFkv1Cdd1XzDtJXjKmmwr/X5DmP5Jj75/CANXyp404cIFukr8gcIN7Wr/z3d6JiHusLFgCcpEA
MoqnF3paK5UTVSehtH+ogoTPU56t+cRIx1MU8B8aV4e3zrjHsFywlM6zd2mJjNMywhSkoxYme0EL
+syD9NmZybKWcPU259scEBnPscMpk5Cj9TwH4u7fd8YKNbs1QHrehaFtq+flLqd9z1rpKd3z/MHK
0eCuskONLIrHbB6RaUo/NxKUuqnMK/qfv3yhsQKF4zU7MnQV+CWqgDAUhYBLBjzdz8n8vlBx0nX8
ggt8dHe1f2H7p2aYR1R5RHHRcA4z6tyq++mY4t851dAbq771Iwvt6Z035XUDLVMgAgRbVGJMrER1
Pfwd0YNVzkK47EDNGiuNyhumnpwtztTKUWCq4bB6fsiiGMfFVrHVHn9Bq6ATF9E/asaU66nG/CS0
+TqrLQoSfPC0RWItZV6drpYmI2ivS3akuIvXHd5e51b/y/HOPExVXgKEYTd0aU/nYiEXcrl2dIlj
AHp9qrHzkjWtzs3Hot8mCnn1hTByC2nuBDXxzc14U2PMfkmepw/WBxdWTOhidCO7Di1BGsyUdi7S
1dAExUJg4GDkUOUOKdL/gM4JmHWO1dw0pbfkGiHvKTce/WumLQCz/gdPKzrk/0T6OjRsLSP0tCy2
G4GHvIquggGjvPeURHQwfSyJ00bYL7ZCn6bJMwQkhSFah6ctCQGtevzb2e+fGl0x1FbPGOahcejH
52qX7kJVHR5kLn8LrC0DVr50xcJSm02XNzzrSW6T6wChGEjLbi9t/eXig1TgrjG8oRLmegUpRmxJ
GUc1/yCwNXsdLu+XeEwBO0YIuDZUh0HS1o8mMAsXuVEo8mZImGT54eX5mgUl+Cu6An/gzQJZk7Qx
LfyA5v5gPPJp2a2f94Slq561+3OA15zc3pUPm3gu6Tmf1yMxiwif5kRAZrp+Q7RrKsT+7yNRdWLF
NmbJQJBRKRo5WqAD65+pcWIC4GKoZELFcDrX2DgRceZEe7NMtQXR2qvKMgklokmIHD/qKaHbFIsG
hZCtaK02s1ubORGAgsvqaInZOQRXqBaLr53om+SosXcuJZI7p4c6NpP8PCRBVgoc4R6qvUPfds2Z
6+7H1S5LnuR8FJSzp3c0kP1kIGoX8Ek97QbJSXayzSVnzpgYixNmtHVnLZyH8SPYY3joH3VydY9B
L6ks7RZtKKllDQHBcGCxizU7s6WEv4CTgXeCVZoRcl/qwmVCGqoiCBBTIScM9aLeY770QZqWFytj
V9YFoq50Q0jiFpRSoSwY8x/TtC/sIeE8q5SbQtAhIMTICeLfrTGSGLSfSM1PE87oj6OuXhyuEV7R
BNU2vQT55uqBK48Emr0DfB4sZOJ5zAEuLKbGGstIfuWGgpUVUPpipSkDyKnfhj23kL+vbHx3ifm8
IjiQQYKCojmZRz8zSXe0NbGKacF5qrHgk6J/of1aEGkApVChzg1bM7eU4PmSXxz2d0uhiN3OTA7N
kwT1ak39QiXBxIpoGnte7X9wmRardwEyWmbmjd+LYmQ1JQD0wz68e4q/7HJ+eWd3f4FlTgCplfop
x/Gxbmq1WPN29P6GhMJfCkRfPzPMIMi6BMQS5soBiB+XEUXv97gcMTPpEgwMXgJYepqB+QMaxb1i
jtmV6qnbps5utQyYrz+2jZpGGUkZuwzdsDtF4e+poWYp93i9v0EInwKa9wlw8fFYT59eejNZxY+u
wQd/s9rkHZprMaMyqsJy1ek2HU1uFlKav+pyjnbMdDOLhi4MgQEedRBQQ/kxkpPhJ6UZgfmq/mIa
h7XZJz584NRqUqFko6q0NUpur2ZtYfhLEoP4NkteQcI7esM2Kkc4PyvGjc3TMuDgo3oT6wH+kjA8
3edw9iqj3dwLO4GXEnMyROIqZjiWEnoVGdvxfijsEicjy5jqW2PEBurkTgaSnC7Q64pZB3mEQk10
m0CRKtrqneVGP+HFL9Xg/azF/P4ECWoB4zglSfT9ZGSYs+RYgRfCYawmVFmCYLzC62Bju9GLn/gN
MQ1L4G1konTTqrmZtzmZSF5NbieN9NuyzqUts1iCSbUsoa0BUoLBirdCW3FejQ2gjgDr1jdng59u
6Pmiya2DZZO5JU6p82oqNVCvVj3tSkhMYjTeCyFdThNGgsKRVF7EPj1UhTZxxXxkhCSkDqvllH9E
lYybU9UODADs5dJfpHmaPIJDAFg6POc6CszvA6iEFsvhGtgXtvwoJeZ2pDlBu2JT8RPpgqH2gOhi
nSHY0DgKbw4TmmN2OxLVM4/Oi2oOOYBEsCmAY2Z7Wz2hYM+dIzM7hsQyeDhAlo2lig24Sn6Z/L4d
3OqVlkcsqIS4LFfux3GHVPU8WW5TRe+rmD2oLMFB8Ht0Gl4hQaI853Kvd1cP8qJU/0ax8y3pdPeb
tJAKfoSGVF2YZ8z0EeenvjJLqhHJ5pcIxbH+KnsDnmDcLGe3pIaSaj8R+QIQCPfKABc7Y0NyJDaM
Y/e/B7ThT0FmH6hVGlKWFdeY4emcZJ6RhMvjReoPyNHNYixJIfszuFZiB0fmqVTHioK5YnDvR0XJ
JS38zr+tS+OTrjOfj1LWEFkS7qlTfoiblbk0RY8yerky2b6scdFKdRFTgO/durzTBy7jmjdInLDF
uAz2GN3glwPMKE5TFWPDGF6t5A6xH6/RrnG1Ofho09msD1rYuA604jBbqmZISO2wM2G8MYR+rrcX
83OmYCblyrSjcloDPm3zsphuwCiJytDYgxZsjD7z+ZcpkzXaC8Af9IxjpbNmO5E9UxLX2aoXovLe
D5e3bMiwd0FdaBe+my20jW2mKEWjffeGteLjEC+knc0Lj/mwCrfPB0fdR7UpMX91AmQqT3Mparti
8hocfqKr/6TVFmWKVfVN7Nunx3T1Gep35r4fc8LL9wx6SiLs+7ugcOSFi4Q3VgSAFVSR81VR8zNJ
BlL9OnFcFG67DmJXgzjAOILMzHM8VQOatavCxiw86kXBPpFYadkQH8LmZWNdfFme4nB0LAiDW5yl
1+MkulZBn65LCjEvfSLw9sQ4jD6WNAIy2NVZKraG322LWSUoC5oNDRdbuLb6yqvVkETk+3PFpVJq
fUJxDSQGqOhP0nQI14+SHEsugMPx5IIR7X27fmNa22ZLTyOOg5Y93uDaw91jzTt3p0HSfxMnc1FF
syRBJVzVBYYsdwL4QDyLtdWhMcaKOP4Fv/dVM+0oMSGmKYS6pqHPCs5yzpF/5HywLmfDD6KO2aWn
sTlddm+Csu24oDMmWmkerRFCwmfk6WvjcqOhKleZw7zjG0Sk98OytF/rRCKQNc0cVkuhgv4DXEhM
mAMKv0PYGD/XqC0X0KwBfgigHDj49zq+S53YT+G782zdTVfjgmxrVZPxW3e401/vrnjxTFJj1iXh
46ZUuJZyBc8WvkVbP2t5MkuAPNbMUTzDjJJjB5cx1ExKb0AKiA3/uGS8vEghl2Vq9HHf4AG60KTx
a91+KvE53xxlVSnmIMI/UZ2EIHNKO3AfoY63bTrjtvQ2q+yjH+0G8/bzxAh329aTcpg41mmvPUAR
IeIgptHMlGqlZGWbQJEm2/cF6RuCoDOs/22tgORx48oTbgFOYMxx33Dxy55d2eW84T9ISsEkN/uC
c2euAJll9oXf6aN8aDwae/vDaIVoMF1TBFkMW9UGX9RI3/6Hzd8rH5VZnUSEWLiT2hVclo36I7gT
xzku3TKCjQjLFV5nk3acjBolx9TsZfiwYXADaFo1WDyDD8Cl7b0TYr4Tj2L8mMhjlNCCKrNgjDlJ
mPlHku1sAlvHyXPHPUlc1kCRE6nBsSmjMi5kQYwL1AcwDn6kYEviq/MS4tZCYr8cWmaZZVkq+PU+
z+jSm9QZg/H5wsGhdnX525asOVdmf5PHWo/WhoH1DAn/ZBEuZAtuaEkI+rV7i9m9ozlFtu/Nfqqg
jcWfAIvLwYRbccN/R9EVw4jTKFs9nwV51BZiM8+XC3uwv1N8PDKmh8Eh4RNMnO9v2SkTv7aTAhvt
CJaoE8egaPW8WOcpJaQhP+W/Pkg+cbjaHvQQ3tsT4BwjRH2HoKh/ueiAuRrbG1mLvesmAZFQTN9E
n6xRuLedcoAo54IHmnIXOX9u5PSSOQzksBTdCpreqbOpwyDRQV+ku4S5lQih87LE/mNWdyaClcX+
TSQ+Vlqc4ASbmfhhnDOTb6LAFsVCOGywUyJX6mfpY7fv+2K0Ry29gWPj53Zh0T5LF0jJrS3GZWhw
VWB4qkb4cwk3GRRSPcN52H9nUfhCqj7Qw670qngHu/FT6EoAlqRnKi2g2b2DOeBl7ea0N1sxBhJg
18S7QZagfOT3wyWpfzeg5PBF7gbH0Nv3x2mYMRi1iSziN3nPGoTTope4ogyDkQBEvYdEf80ztZIO
fv4+0+GJdX2yReQ6dg7ZTvqNn1r2obL4q7EWNX8HZI+VWa6hANMrxzBX3WzBJyMbDXBYze5Dfyjj
6O+cfjiDGTOQqLIO36XhaeZrnrDtDbk/X0lITrayWIBTOq/TwDo94i5i0p6krWGPWY+047D8ifDN
9AdBJ4sQTHCURay+i07dfq481YYwmB2k6FqszxfyuhEYwARSpagD+NAz9dMX9/C3a4SN3DtE/Teq
nAPmHUeSOBTz87p9K6lLXv4altDa9Fahy3VbJRv/jCoJDoX1kQP/SHSj95iZ0qHeFzbowuCHnYf/
/0I8mz/LUc71vbd0pJc/hlQVhWgDIt5+O8aO2Q4+07uXc5pUNTrZwC5YPe/OkHBSDWRlBH5gBE/L
ATTu1twm7qPkUxpN1NWb3IkvvrIbOg174GmtZf35L3knP7ZJ/aRum4SOOUDIK42NHoQ8D5kt3NTi
QGURGqSdJTOUbw069u5460Zz4nKQVR1l0WI/fiQP01suW8DrnIgzWHIrG/zVACppSOCceOqDdtMa
04F8g7kq7kQlQUc9jUvqyuUlkaOxWBycnt2DmtN+yO0h6RLg9cdAF5MO0bQIv/0Cd0Qcz9XXnIDp
mEhPYY24FR8mBb7c31cdHou44IqcIIPa8WNAq95VH90ZVAvpafST611bQaW5R+E1MXXNogVWSusJ
Wf3jpUt9pmRRh5/OIC/R+9rrOCpWda6YhtfaBGYtGxX23gEhfj9xCrn2JLA04vShIfK52UHSmyek
ec0zHbTTobyefmRBVHHqCz/tErn46k8G8OiuNNeVzoiNbaiBweVORrlOd7yB1fRxo3zxkPSTxaWz
Bx2x39eDeeCnGgPLdcjtbN1B+CGp6meeij5RNIYyiPNld6CZsqTe15rNOKbWSP94wGhknOP9S4Ni
GBibCG/8SNHfqsGfNBJF6aunxK1usZMWO68SWwu3b2eOFP1mfqM2ftMvcl0ah2TxoH948WnJ/nMx
6E//7cRSa6cW7Bx72u6ErrkzSJdQZ19E3wbx+erGc7HiXyQVUb3pOChHnPecJm4p1NIL0EyTWuyp
gtDDMsJwoyGAmSzlbJwEZSC+oaCQ5Qmn3RmblGjaLrkT2GZyiCIz/9Pbd3wDI/LT8MpOR4F2AhWY
+8KW2I8S5/4eubBldYkOTAT+IbMBmJZ/NAbIXMR1bgS5Lr/vV88GECrGfiJFfAdFDfHxbI/BiHKx
JYypaqZZ4fCQuuwBPh9RWURnctIcK9F1dMoVSmiIPDVWSmPZQRSbTYvdmda1hC8tivkQn8H2Fcwi
rcV37EiBjLfVSZ2Isywy8jnbp4hiC5gV3gLbs/nqqRKeoG3g2jSMKFhFcp6LqzJ5Yuwzslh+uwO4
RjZruYMH7CekCr/cR9/IqSE28anxP6bwSuoudKc1/z2soOXxhYlCZsqhQgp6jZbjXzPSgppJQs+B
+IqSKGq89gyfBHTjj3QpUHCifYW01rQBeAoo0wtYIWO359CWnWScFh7xRqMp5m2Gub4Yjs8M2OOS
JYo7TVVOG8FXLREUQOIDmxtPx3FVuhp6jzF6UT27VJh3k9+M1WfNxkob50aPQD1z9FV9/FOJuwnh
zeIcKdUPrsKSdQodtLIRg10WHiQPbksa9qDR5u9MIHSsVPmUguc8DBOARQK7ql1lPpjI16grIDN2
rN3NmadH+8l/H5pJl1SnIbbRRwEEDkEueFmsX/kBeqa6LvkOwUybuDxns1/9wXCB9QTP0ExxL2WR
KfDwm4hrB+XeZtwBp4n/kWzp4r6Epyjr9Gx5sM/pTIXqHnZiIzXlm0G05qiM+48G6DNtESAlBj1c
w69inhQM7G4Z4Y/Jimd69rSnODZNQaCT9F8ztryZFSzFv0KnE4ICJBS1gsB8KLlbhZA11oEoYamG
q/wQRKzNnB/5OjAlau8agiVbYupx/iXgTc8l7rwnVe8vDD+TwBIvF0zYPf1S8HnbYeJO/c5Mb3sU
akYc4zYLj0wnCpGttfm6NX6RTUlQ/fgGvVXEVjPCGwhvbr1nQ/KYYVEzoUIbQe3flu6Qs7HT/nzY
wzD8E6nR/cNT11/Nh/z27U2Na26ipeuUJ3ak/fryDZNliKq1ENJ3EHWnjMgYC0S2nRQRUyC9RrNZ
j/P9lbME12UnK1q0JG/c2iTzOtvy7sjpxxSRkmVrdh4VGEMKRWgVejNkiiXHnxa7ffBs8JoHMqmr
Q+gk12JVf1XhbfKYdK4cvL23tzPmYazW7CB6E72DEpf64/QaoJzB8oO0TPNhtC6UxTmbGfIZSBWq
AAahLMZ4MqjnrysH2A2aLbsBqxitTbbV92zIW5ocBzt1ImZRtkxz2IRXyUAIpmP+bonlhQhB22Jx
p1VskFxJY9MS7k2l5VTx4/1dSoG5l5B0KGyABEMsP0oqxVfMlofSBIhhj54SVqOo03co+JUX9jPb
wfULBv1LLLU6Tm0mfUkawQVq6BbAVJIwJduJHbyw6wdhlTlZGV0kuBtHwEIALTuaJOpxSt3B1Rz4
+qfzFlraW9cyJ0tC4hE8gWrp2QmcGNVdiwC6iXLohEJLfBq+CjnEFSp2NVRlz+M5hvFAE5JKn1gY
4kpTs0y35fn5yDwgGICx9/J26iM+KUCZXR7AX/i4AzTHj915guI7oWOyjE8469P7KS6mbeWypYCS
OqYoPYcRhcpFmfgls70fWSMTXQWL4W6c1uZU1GFHA/PBEi8DOSmDyU3lGsa6Clc1rHOyMEAGrBgc
SpHZ+ZD449EplYJlI/c17rKCAqMOko0HAgFu3QfBajWD+c+LYNpy7VcVexoLM2BM8g8HTdUkD2yR
v6VWWV2O9fxhBQXkj3m3c9EaRgMXTtBh8r2qmPo+4oiRzhJ9bfvfrrDe/jXMy13uPV59ot5dV8ya
i60irxjsBK5CG8QhT4chBNWqsRaIqFWdZ1DV8AMtxMntWKcdIZpAfVzSKZ7vKg5qGSyAxk8XWBry
rQoBMPIF+N4oagpugGm8o7w2GgC9e/aoB1d81V8YDd0kBN8MIq8knO4sorBpbKSF2FDWbNYLyrAd
zwtEmnvHYhtoXybHmyJXQanpJV1Q5p3Bjnd4UYH6UUNwa73IPrKV/VdbdF0SrDl6LOhYZ4aKyLYy
8RWG3KqGdwPZ2XyBGiye9rZblS81alvgpL3WIVL2VxoZJEWZMKGDaFHz5R4CrymsF1is9e57T5T1
ioveNU4Gc/sgUR7gctPUsGBJZF5TdGTYO9q/riJKYgFwkxV7A7hpz8A7lqJnQ8ZI8St9n3bMgYRN
ajGP++UyDghjwCam8xJjH4Cc8dv/36/A1/1ClQaCQoo2DNQDsugsQOsJ1AFmjRhjhIqF2XzfyQKY
BdSRMpb4gfqqJreaVmGNBCGsYD0E6HHUTzcvGKi1EnHdIrXuEpvPOj19RlRAyWNMHIEqRXiiIzQn
jtK/7Cs56WCcflHPTOpo4rwMyGeacfzXd/9ivJ/t+B6mJOQk1cyMqe2a+In9Z84/t/1r0bi5M79H
1REVaHWr4OTe1Ayo5+vG2zEPDyPZ/u9LpHRE8WdUbal5O8LM5C4X5tigz8l5J/AXL8viQjVedX0w
/SPmwjxgOfJ081UtUMJB4aTVrTlEbWCDVmgPPMAXrDrxcS5B5S5rLClPahmutcdAzgkdz7H5FMHP
Vaqi8K4uGINDl0Q7i03I+4PvwFyEIEb3xqo8kbRkGRLeHoNJhg02HoNQ4nOK9VYuZZ767Brc9S/v
2jqCRG9RwnjWPQQvJMFlbOq5pKp1jLPkFRDfWqT1yCLZVb2/vPXsIPO7fU0GdG4Ojgkz0hg1tTJj
CLzmatzyv2bxdTJ/1N4hOqI4dsu5VfxTxXVXBMAbjmwGW4GeQM7CvHZc7IK0BFnFddyoUQ+uzpCe
SDCxfcXbf99Ss0R7kw7dtZ0gLJzrzcAc/9cxa24RyOwFpyVH0EcVPdNyvZIPKU2OoPQREoLffAQp
QTX9qJ0FCNx/PkktcqmpLq/qRDkDXDanyIW/hTPiSKv92EuYo7tSxULVzD6SRWFEQXZnKJOW5b3c
C1Gu0DaQtO5fM4xQyKzATN2PZ85VLJWCQvkoZwXawhKyqLTYdUTMCwH68c44ByxkpAFcY0fY27s9
xQBomhz3VdSoLpcRhqkrDurZV/+wcRwMhlMYgl6sB6GNLW1cle3/8FBcnHEE6/eyUB7CcnwZTwxt
RbGtappp8+LSY+DDTxXGj+47jBklZpKXHWF6j9ExUQOhuJHgGb+64+h43zNlnCz6Ix1UAu3vqGPR
ucs3uzBEDdCm7n8Kf/QPmDq2uilcQR9TYzRZ6Ic6TTJaO76u4ia3wL3+MYX7m6lHvIBbd8fJg1NZ
f5PHDPcJOvoVI7vOy8xbD4QUmD+31q1zlCqImbM3Zx0ex+UcznHcBiBTCeQjaPKP3iZfmaHTFdt2
gOoiJ+3hRGjnaluIYO+cFvBE6jBHABn0p6diXkyPgr9no/5DvPN5jlVJlmxMPMXgk1CXMxEEI8va
9ASgascWsdwtm+k7DvSPfsmSLmi1vX4OC4HCWMIlKHu0sDZdPolt/3thCEf0QKoxjnkKnqML9oRc
Dh3MrrqpeiM4CSH4H0obJR08O+fKex1HHh1CxrlvPJacej6D+q3YVoZ5FObe+O239HXvPNe5iKFM
ldZrTm4gQoGsgCyKcklO6I4UZa98HX7Ap4N2BojEqhftadiaAD7YnZtYBTGSsru56yYTSUdmZIo6
wHLascrBX7Ma8ZwyZmniFyVgTszui4LSy9aq5l4PKekNUCCVTg8XyN1qkERmq+FTnrM9HByEZWdQ
10tOx6t8xj65qtHfjUmSFptOMqiAhtWH4ivsubom45w/cwTaek1acL487uR8mkZzG/y0uxMHuY79
Rt+fPZlP2YTb+4RgE3yNANfcxTcDqyWVxl5sOhFTjSzRLShmD1IErS9CPV+4j6DpwWjxfL/qmxML
+NeBtT5mDSdrKwKAlGaMYVHfVKS4bR7BpF7O8sNcMQyluiGNEBxOuq7QK32z85mD7LF4PNFwot20
LlDQqmUA6v6zYe6b4aS5hKSRZ7D0jjBvFMmsjQAMOaAw+LmyxwLlOwmMLEC/cZGSmwUUO1SbwI8E
qW3Nc6ChyPZBezXDhaNWlWmPigHvkU/vMi8TjQaszjqg4xxo9kXeSaZZzBKK14Gj0MTFCAUS6Vae
6yEbiTR5DemyeDLb8bU7GE3o6iCcm9D4ARPNv7XQ5xfn3sTcY0B2Z/pDj65UxRHVMCuwRVdFFo+Q
tHYv9BO+50ccJADNw9Ae0CFVR9o9Tv8LomjPTFqhGc6NUEPj8wUrxYirLUJ44y8xtn7QqCk3K/su
zy2KHJcopGBD11iOVXK9ru69qpgGziFqxK4zDtf4wa1yvfh+R6N1A4v5VSGLP96JC7DvOYwpbhb8
et8UYFGztVkOg5sTbIiNVohajz4mB2SY6gNDtYRdLMHuhwJmefOjwhjAPmRtrA5XIuqfd5fZv4OO
MqFcgNR/JMty5IkbXekovsTGdkW7drf7pSP6BuPj3GTG7ZnNO8KzfxajreNENuWg++QOyagNEyMV
Nlg6j1ZMUp+1HI3hRCwiSdfBJBqlcLSwPsAnsYXXa59jBEFGYdO8oR7f0auK6noD4yHvp3mrKvEy
KnIIJqvSwYwxxeN0GHISVM0v0dOR1vFa8PeaMV+Eoc1LfScbz8sMffgD8zWGuGDvbkzEpKkekTLx
9XNoA37du2JApNIcwFdoKqKbUHO4Hky0mudRvLfad05sADCwU7GEf7VFKyKoqtM91Jb5D6x01EjP
s5PVvNWdQBq17a4yv7TcZF3kAm4QTdapTy41fVgr6XkiEbRIqNW7J6NypRN2sNe2/i8SA66sFXNw
l6Fx+AHEvQtlz/Yqfupy9v/cs6jGmEi3dG6qO3xGRcEtSe974cCvB8OSuPMNpHUDVmce9Dj6RW3S
lW8HcOJKyvhYcKMUnrfT8Z1wA8YXLR+fioI6QOXjNM28HgaT095mWspoNvnM2EYrCi3biUofQrth
N6AQc/iPeDkCudHqDj44r4j6d4msysjan3hBfAMoljgBxsfpJGXqbtp/D4wICGXv6N76JSC8RNac
zq3LXHyRyUyvQMLGoDGqQNksPV1FDfvqVZbMUtifyFETPUuxWEIyd/GllguzkS4mVAYfU1rrqde2
4bh7bb5ogpIfwZVA5jqghQtVMLz5EZ7/Ul3+4CzkPPrjvPxYH0DqnrKVCbsVmAbBXQwauVfsEm02
r2hFxn5j1kkUAVHZr6ZMIxtZwWcT+c9vpqvG7JA13qB0QB8tKdYAgUzxgUFNfFOFr/uQGl1dvtfJ
348fq3HkRYx3/bnJVUrLIwJ8CqeM3D3PkuKqHq/conT+o2BxiNiFWiQbzxgXCP0dnla0sB0Cp/5G
kekaDvSMT+aGVByoq9y5RsDIrkz647wHAU8SwL6D+fw5cUzBGe8vYd2z2zTjiovsNsNRPtdsXbJC
//4Qkl8Ewpxr8ArRh6KaH2yFcSvCTEB8UvTcEe72Khb3h9i2iXG7lPPFPMII9jtdWo8AS40QADgJ
yE/f5w+Nvr4oJm1toof2ZEX0tdnn4+L9WB0HWRdvPTLcnpcCfH9PFYjphH1Ofgt+wILv36GXwXn6
mI5vMIyrVZ8hK3lxJCiQqOGCCl/lf9z0j+xc2m3RbUrcfekctVvFirpxn7QLxTApTCw/YUqtCYAk
Lj7zRM6yzCg4MtCriva7n3K8YFM4J1dKRzcOaZOETYeUy1fOSUal3UvYOiB0rs85XAEEGRpXnDj/
I4YEnoPJvnBdKr9Hg5x1neKI6Ki11JR72+HVDtRkyqIkvXwLGaqoHkljJ53ZkhGMJZlyJn196NSP
JLedRgtFqSdIZVb0NdUNGKwr8F7CvYnFz6iiUtTrVKz7fwe4JU3cs4s9Cu1Oyz1AhSiNnBdidUR5
9kABNaUCjBwT2szuav/soGqoW+9O/Qt8mWcH7X2bru+vPaPRhsbq26+SCQtHVVPl3yMnEMjFnwou
pgMwN8DGF1tIPdScN3JEwejckplSSJvB4M9H0DOsi0aU8adS3R61mmNy6M1vCL6M7+/W+vtNl/Q4
XjpqMTncIx6Tf9UbePgJdAxnGHpjVlHWydaVJC9ZB+O8lERQ1rmcQhPH60Qp29sy3873U6m68kZq
Q/lgC1c74FNNuKugqrVGPOEvg7y4zQkKEAHVM+bdxGrn5oPQDA9qAZayzrzzr+qB5jKd3Q+IBqtO
srxxwwhXgr8rCOJNKh3EGsDOGXPXC/ve32v0MhmlrniCgPsn0o25aaf5tX8Wkpv5ilBxEDf8UByy
djXf5Xm5z5yK6wyvbBZeBPkEc14k2GiyBH2i3y9qfcMGluie1aqqm4qX7HGA0/FVoq9PxazLgTKv
YnlpR4APf35HCgslMCvDtTMz6DE7g1UaHtsgoi47hUbkxesFrfxBKV3cgVnDef5H/ln0VSC8QZqk
xDpRFKMdiy3PlS7isirmlo90cRTqmnxAYm8plqQJ0TKdY2Dk7omhxtIW/eHXXzkg4xvP4EZJvbH3
3x2FffeUHglUsrMwfd1i+Rf14gpGbKK7i/Qqe5rOuA/qbEZs8PHIAk0NKT209NMinaevyohQkJUC
tFzd0vZby7sS48/lijmWBtD5FWNEjhu7z7zPlx1c2WkBVyE4DUjVjJQCxKR6tQucJTkRlaXeM3ee
8YNprxSUdbyuRlNXslhsx9xb4BxBs4sUY6jLOg+H6MSWZFJwCOEEKzcXBOCNAdSSn+GWqBOroYM2
nU53WsgSHUgMPTIdVkHFYAyLpry8e6SV3w5md/qeZ50AXP6DdWt66j2xWx3gDcJBBhwf8yXy75ot
Trg94jUSnJ8l3xZ++96M7uaX/oZa5BYsO+IrZsDn0/OS9Q1v8I3Opd2xEtmJK500LG5L+dKsa/Xn
cst1tjcsfOZZ0wFOrbC7qDLY/yPN7EUrYvCI4lKNo03LVqJpPy6NGlYXjeKhFB/lLsb0bjwtfK/i
SMf0xso8RcY2ddY937BDuPYYH3x2SlUQwoGc340c5YfAUzL/OxSCH/UiijiZ7b5w+jmCisR40ugr
e6rzjbpm6ZI54lrf46XVPdSBy/RN4sIRtuIGl/ZGWdN0bYPB0q3264C8vQJLY2JPqWNCaSp/3Bng
T5ItZcHR/eLzGG0mt5gdETTlAJ0oGH23/KE7dTRRjKIASgk1JhBhzg7AEdmMlkCLnzorgDRuAtcx
Fyu52BrS9UACgYSI4yEz+mRmEUYP3JgVZLTqZNGuvrvtXpbSk8Gl6ivy1Vv/Cb3FwgN3OsW5qnTH
JG6czhEnzgmVse0tDC2GVtZKcCdcVnfXynYEykFtKC8jWHw9B2uj0QXEzX/aowC1Bst8bLhtIqek
fgeTerRXAhj2e1ufU1ta0HjmNc5L34Q0dtnZb1MBHtgfYq+r2DQnmAe0y4VsQ9e9jMDPJzM9TcGf
ilFhBXBcHqvqNG7OHtce4SuW3b9Ak8Tj5hPzTTP42/NvDU9KgEDlDhYUiV1SvjJ3UWNuxwocrkFh
T8TOXEWvzVg/SIx6vykutTBzHUQbwNuYXd/RYjxU5nw9F+I38B1/ya0WiSBU0UwL7jk7gVV7Pch3
Nu1FK8ILXLHrWVmoPh6H3xtpOZ+MpDaXy8maCdRyuogF8BG4qjZBuov5Kj25o7BgyIeXI082Gxro
JTdsg8del4cVPGLu6WI588MiXHFgyxSEh1nq+1mAlYfNRsxaxOEVsvMFNDLp/TJQWV6WAcMmBIqh
E/Y0/xWHxkg+Xx3Su4R1M4vyM9AcxI9v+rRyaSPrXZI5ZbjIIylwlLfikl6hkyflT8dPziGT+/o7
rIEfm2dxgdIS8WTXTuXQGY+MEv2Z1cQEfxZ75OfC7Ja894RTRgfU7Td4RWIxZ/7vMWVqn5CwJWSj
wTq34bgnJRDZSc++QKYgz39eh5R0c1jLeA/VfY7KxMToY0fqn9GYnSo/B9WaZL9I473mnRTycWQT
a5MI7hZxL4K0UaT0V5NdMghy0quwGr4bovPDmuX2Ce2FT5wBwdJ5V2Rp8ltn+WdDlgQ1anaiQNap
BZXYNdkbH9LperUwELidnW12R8Puyy8iwgFIfkr9+Ig1KZi3LqLtmaEimS2FtCGIlrQp5+RIyXMU
RANMoxB1ae8o6urVSRJqgXNCV9hGRmVc6GcLX02SMPe4jFr7QSZ2D9PnGmCmqPbWbqH0ho4RglRf
lajbNxpq23nQ94M7dRYy8gudXxX/dLMIeRprzApG8fh3r3P1Klq+u35p1oYHF9YkTV24LZ9wsmnV
bdEZqGKwCvX1nHwH2+6z+pZt898DSG+J0O05ogTV6Wao+4PbLZnLYt0LzVrFgU6I/9m8V9sDTgLD
WpZHIbUz2qzQh+HKp69JgRVDKz14mqLyOGWCc0NmD+l/atSbSKYhBmcowiOG+P1Bj1FftuAMwmyL
vqI+enVVXMqqLo7ToGl3CEzs7KPn6yv2ezG4PDskOdaX7MXzoMo2RSrHfwo/U5hESPp2IJiqGZGo
bo0sV5Qb3eFgmlnHeDh8oydl87zHqThYGQhn8WI4I04lVskkl49YBNDR8tE1bB7G6rJ7JnfUGvpJ
a7L6I7NUhtQ0wcA+dekGrUYYlCGLdsSirdv2w2LGYn85sBx2VgoKUeF6Zjpa6UpWxj/TpMS1lDpA
osG8IMUmKHatwnPG3asSO9tj4I+vN4rYl+i/DHs5FcLIwjvxk3VGLQYeWluds676OIpR4Mlq0+0L
NWpGp3gkvDEgILEwYSf3rTn96ui51Hoi2jWb4F33Ey205NoJDfTJHI2HQR4s+Y1Ue4lwLTmMo8i5
UNXURjEH15+eUa0r8mVDjVR6noq6bpf89vrD7uc6Y/wPu7H9k6yndpJlLwXqABtvMqc/Rg/uIlC+
5cWDL32iV5CfdzwvGzsslZV4lpa4GbKKFtbqtQ6MyiGRMl1y/H7o5vXzWR5+W6EoFfMO+ujt7TXL
8tQ+FI82q2Y00JgMBEp3kw/VmrXp2mNTcXEfODLUg2ZrbcKiTk3ZCQZve0t8vF25fDo9zPm9DKjq
J9wya1J1uuHFDTOsZSc5hOPcnhf/rkPSKfiYXb3G6SAoNT7D7lbf5QZit3kDSZrokdGuH70jWHsC
4GAYsdgdQ/XrONmFb/bck+au6mRX+u6vBkcOxj1vvKaPjE5ROHeoQ+TzfE8h54XW2DUr7jpO4pJS
ApqrdlFrR0rfwfy9WaOHyycbN69qnTXdO1a0d7DVuoFuosMI4QGlBlsma2brT0cPCEYIhG0HgZ56
q88STxc6dgWe7TxAlV926FKOMxk5nJSjp7ZyUkaKVFWrViCWhRo1cBM8SoGe8iIwBWhEcXufXruB
omsS/Wg10CVWRVNHh9pGiXDUqcOoiM7REDbTxzRC8m2XkszAEjnmLzooumV8GBes8z5/Bd1ExPvp
OnuY5rHG0eN/T3OC2NgzaxMsyF1n49OFVP2jSH4BF9gwE5UVtmLE/gggJcl5rVqwbNUILD8emque
VgETQ+UsApSnjW5k7s2Hrw+FFYmx+araGpP9BFYhwV90FaxqrN8dn+I/nZVVyOgw1/yhJSvf24+Q
YsSPgyh77UPXrcrUQifldVY0y6ZQobfc9psAggCKfd8xM3Ddc4jGp8TQwPeF8ni885soHsAqooW/
O0fuCFMmTRx/SgjfUs9ulMLCabP0zYGJnW1N0oaYeeecnx1jS+Vym/VdWHYXZkkbPXz8LNkQ6psT
NSKR1ixrmF7m/Wso9g43RvxwPOS6xVprt6vc5tFhKYdKFRBFR+GeaJ9dgyW4dBqr0WEr8CUqJl7c
/KRo4azjcmoJ+Q0Jkxqr+6X6SvBlpa9AYX9od1HnsMCWJVnyrze+3SHuvGJopY/XhNrICB0ocsbF
mGj+1A1bcymRcav5OhVboH9eUiwZSVQcU11avZAefHOEAC9gKFjyA9gwuFhjuaTza7CqJcp9PnI2
RLFak+PUpaBfDCPbROtyT3wX+yTHK+JFcPwch8SyL4C6eEEE5nPh4myNqGp7WYZz47Xfu1/rkZ35
7Vx3dMBvtQ8wG+yuOSaYI2KbkdG0nKrD6V6Oam/9BBFtepccyTB1EfyRia2hcuHydmt0AYSzftkm
6r02tV+wSeGDEpCeUGHEgPw9RgO+SdO4HCOLiCyWgAp1attcc32htQfBq7qno+k37btLtTeAxzY3
8Nf4OJM+iNqF5gRSHYDrn8SOh57LTecpHNOUzAgdtMlVpHGDT3x3L2r2AUbxswxYeAnO1oxh7kE/
tILi1Eeh2hswAQPiK/3vUpsSYki67q2LQ+gVWBiWKh4Ehk+0FFSKr3gICpMSA+6ZNapzblXoikFI
yxsMFOi5KIfz5SR73vPFcC7BCVzGbIxiO0SpkBMAyZbJQ1sAFc/P91hqEfgKcbAaVZKTo1/7EoWZ
h08LfFd54xKq4OGREfS3zswFHREvAoAhxCjfD37rX4mZ253chRKAYuA/jDqHinXexpo45dQpc2Pd
St5Kt/LhDvPNtRN1SWSaEQ3arVOOr9NqU/rs+JIqQM+ux+tahtaySjolkvN8GYxg6tMmLSh8DI9O
PILQtR2T3kBLT9ppwVDWPPDRJi7bujhskwpvUB0IKBLmQN64tvwjjE3Rd1hwMsY3Ojrs9esDM0J6
kLYKfitbhWYTRV+GgtHBzUkrkHoV3EJLDSz0XvgzTmWRqTz8nZ68NoLSGN+vs/XsbVYMIIPjdNIw
H1bf17QvEZ6Og/tYmfwflMhHzORfSo6c1qzsp2zNbQB/++7M0rFX5Q8GKF8du89zHaaJzvB/F8a+
f4cGbzO3sUuryDHdtFmJsMXTCQNy3rXuGnMZ2YteVw/a2DGO7/jAjlT7rwoTS9EsB6xFYtYwQZ2A
qTo23DRHBvoEFEQmtRe2NfIN8ohPJ6trY6JnRrpxL5sdsNCDQ4xkrK2yFxdH0wDlEyoRE0Osmuon
wPgOGZbBX8cAr4+ZVFtOtRGVi/TXjQVNr6L9OH7N5GPO5UnrZWWzwQ69rAO/oOM/1/VaVRobkY1D
nVoF9fEfjc6+B9z/dKwu5aGXCiUtKZppKDNMt8R2VVIJI8hnfwxWHpgBKGuvN1VkU/8hI+dmHykN
rR07W3uJKESjFmo15skWOGdSBjsEjSjHNa45lxSAyII7ITUSzawO6T4cwptmgmDwRojbNHH2S3RY
kskFrsi6y7fswZdVRUB59rQaLGBJ9W+MyqQ3WAgz3edZYJ8LQ4MWtPTm3e3k7TWKAr6Aw3tAfesy
x9p6YHxs+8YjvzQvuBRhE+lW4u7g4N14MsRoM5oQjrNQUDOeH4LKB5hxjgb+JlWEtXKT5j5YA4TA
1PSluxv6BqNCj8KX8OxKgnF1qFgrGXsbOUXXL74H0KLTVwXRrTMcv75OblGmJBcS/VaIyNRaXEtz
E+bQFwTWTE/RGC2FqWj74bKKMkVBdwgdcIAnL6dK9AsRpGXZMgSA28wE2IsZQqH449+DMkDjBRSx
vgEVpahTd0dBNsjRsAtUaBzmjkzTi0uVq+nha8cWFsXxDtMsAJ0RresI9G6ro6gTrol9TxYnidsd
WBcR8UM6Kegfygk+Sp2v17AUkW0TWHExLcw6daegvEs3RLGqA0QiLcZw2zcFAd5mKcaUcTtWbEdS
tf4+3Y6D6CEsbZSWccHEfp0Qjta5KEFINywZ+2hQYxlkw7134JcxzT00qpbYLBzsBGrw8pjj/6nF
xvWC7+YIw32fcXLP6mZpSJx5mxKM58rwAnZkBs4suUdwlCS/9RO5xXXoYu0pbbuPJ8alUvconG3z
enRPcJvP3MUFhhTjsOe+8tdWzCecfPXHR9+3nhWPMJgmRfCuYYyri1f4DUHE64FdvHF/O4/1PZeu
QKtbjnEknHE51cFbkhympF1i21qZ3rqsoknfzq8SgYA8VRekXaNxL9Z69mR5edHVRPK4UWRqKe23
PvBRth7/X+B3P0+nw9EJBF9lIsIoduv1BM1yU2hpqKUuYmmguMhSh77P1PzoM0AOiFN3HZf6AQ6i
w5JhZ6lHgrdHdDJM/r8gHfwb9FRsUSdsdQtB2w0hGpMWfOJ7C3UvWNGlspgR01DS+waIDjPtZGJc
ASBykUDDOocKzCYW8QAw7ZIl4xUEejQNFsmm7kSBe3y/rJLix2wSO6j3xzDRIkfCaj/jSyn23GNP
/NF0u7ojjLwH4+UK/mj7DptaiTxtpHTiqgZnsKOMzsWPcp4qJ29WxZxcMsM2UwH+3VBgBgxypiRK
VRy1ua8+YngfJ+5nY4FbMcjaScbjHg/BSEGDyl/Bq2XILR+4wSEuA1ADthauNHpM3vQnfJMa4iJ4
9okVtq0JCvPFn0bzGGPTXOQYaAxqb3cDyaAqNFrC/bZy4WspAMKGaKfznUev2KJV96PIKTBdoTW+
gC1TWzSIcQkZmOCvpVnvUyBsWZY8QozUpBUv79ZTvF5ADaBAvdoO19DgSGblhGAD8dI0/m3vpTKQ
1THKB+DI/z7pxPkMD9bNlr/JOguLucPKM9TY1I6zcGioxzXHeoLdm5qkTFScSXZcC84bk0HKBqOj
SLKxLZeImdI0UvFq2RD7JU4fDSfoibWTParmVf7bMM03FXIa9sLe2HxE1SriEwSThszk4uGnECzE
6DXGc55/7AJxK9AJ3F37Zq9OpaIEI1kb14oh6QgK/JhReB64EJ1N+e0sTCX68INjS39HaXc9Fw/V
zHA+igRypl9aFaCda1SrLl2jRjSQ4TQt6gjQHFnxm0O3xgK+t6qC/iPFjJ86m8hGp5HirJtccuFo
g0ACvm6SbiT50q2dJkvN9mQ+FxdtX93eHI9f/fFHc23XWgAtoC4L+MqKJfAueDYCKcvwUZlsRBn9
a9vSRffH4fxEb1OOTfCpJqJbndIBZICJZfoveKekvkAAD2f8DvNaJ0SB/SvuFiD6FbEGGR3QQm61
18YVXm0PmMkSSqaptNRXz/IoE7xiZuuIkwy7mh0E/Acgfnt5EW0FLCqv5zmsLNXH+gjCIfkjzl/h
IOI+4WuILg47l7hg1QwNIGMmJJwtTWopDP6v/wuUVCiv4iTYDxODfxu3NxQjE3oA5pGFAJhkDG9z
vweJPFML9LedbEra7i+jWM68ncXbjqnti1wgjHKlBKEi+viSUsoS9wBPhNbMxoytF8M8BeKXs4Jx
oYXJ1c0VXjDUK0lLcyFFbBpfFXKxdodixACzRo1GG72t+iBq3fIEtfrHo84H9u2pVLvQ+zxjb6Ei
aB5ZEQM/RgeiMU+bk+ObX/Kt3DsyHOjWpzNReJzlBnJbv34hzhq9BmuNXrNXM8GAyb4esHPjNlex
bfijXR3vrmU2fc8nDwUsEKWQAnV3UExYX+0wPlzSNje9wwXsnNa9jw5ESk+KFdgmPEr/xDpXljvF
tpvNm5MFWyvJIMiwX328CiRRder0jZgg/E+jac9ahOmS1DjYYIULL7LfNk+qWaDQQQEprsToV5xr
nznPofpxIiGRmsL5B2gUblENgqvQBAxNhEFjCaBjuHdFusWwtuleSzx40apHgrxKzqqxm2xabNie
dPHFFV/7CUfrZ3y/e1ltPx1uPfPtFx1l40qZoQowLR5PNeFaMDzxen7ez1+0SqV85duQxOfftum3
oofpCbyjnVduG+AevqY62rlz4wCXlrNdl+aJIhOB/gOxcpT78AjPAmOE4FZKuwzg6nBecdZxlons
w586zS35S9PcAO4aul9cPLpXm5ZWbdmeOQN/baIKtZUec5/BXf/BXlGEhXOAxM99xeQZCmDC5Zf4
4RVfQhKjY03IS1T5EsmuhYwJTtxubw2c/k2+CWdBJJV3Cox0K2jMzF7NRhPI4/5khFCbcU5HyYJa
sMzBiddk6qQxzkCWuQmFaQ0Vxz78yvvWVDyihGS8Hd6IUgOwROEjSMBqg1Ms8+ZjK66EDpdllp1o
jeJirZzLaPRg+5lWhkIAsGWRzbvE53ReqYvbcFfC6wNEDx1h5DE1nPlCzpUKCmO52WNbg4aknOBr
o7oUimLk1fGmyLXq8fLZg0yfw9j/555lG7lfkqWp0mdBHE2L+7RhXgyY3UmaIPnybLfAdTIQPtd2
Sy5Ly12tLrkuRYluk3URHDn92amrAI8GkEFL89kC/Fv5MBIOHApyzu6sW7bauRfbfEUpE/T1RxPM
BFprOmssuBjdYjFxCfyavLYM77dWJVR5eNchAUgfzCZFeOQmCB/ZAl81vL04pFq+/cEy+wKH4/EM
80OSS/ZyK0euE1knkqu0tEtSNQeXLfZSqlFlLO3rvfo9v05PSLprNYt0MSLOA4ugY8E+/py+YYPk
6ZgK1ev0WpZBDh8b6+HhmeLS8duXamd3VQSwJkTtkc5gbkPdzydk9VoL1e/pV8rJOH5jSph5pagh
PrW2U/BBSAPTN0swSZdEAg74wboILIxAye6TnX90eiJGRzBWlCF1lZR1C3r0D5QESOQlMhmkiJeA
iMmVWD+DrNof7pbnCkOhQBJdfV/WwbqNv6Wv5IFtbpZy6946wCXcjsSBrH4ABVRVMIHcF3SQoXW9
zOnjNskX4fpoxPehpA/wqvEYlExUr2QiCGu5b7paUlk/BXjxeBe/XFI0fBLosHFUD4EP8xz6PYNb
scCM9fszYcvNfSj8ER2+2uxq34twYojcUXrntHz5SMEu2jNUix0jYf+vQs8ZzIKhv2ljEmtTxCwL
De5azu5RNm4wbYinZm1j1kkX3aYBUFlDWLg49d84FHUsHDYNNKsh9itMSzo0KqpWLA7cUvwD/fmD
LMO35bz6Dq4JJVw+Vr41B9SGa0FnGYIykhtZNFrTrMxkEtolPDpvZrDVAwj0BSLz4K0G1i0Lbdb2
jumD4wmXIOlWUAGJhnE5Tzoc6EZPUU+YNmiXFcfmUT5WlH7Gn8Lp3v2aNFp0nhuoRGMVmDKt2ayC
Lov9bEH4Wivq5ypnp7xvvX+KuzCmMCNZtncWe8TZ9DhPzhmHof/oyvZ2xNB0iRjLV1O/LJjbnn/g
cSpzTUMH5He+hpvxQRgbH9EkcmuCptdtJhdLp8k/0/zZhEwLQWja9fkFN2afbTBH4u6bm2bW07pL
CEMHsKBW+5SU++FqaEQVilRp9HDWIMVdgldVOiq28GZi9LZTA20Jni01qAWp50oDYAqDDFDarQMs
B1N0TBn7Br3mPYAKbNbqQ2GoH6Du8lw7kBWfay3h64JyccukzDhvf4Xt7gY2cVEBKFA/wP7TkDO8
iqJfq83hnb6Z4SoEVl+t1K58N/PaBUmrMDksB+T+z0Bzjo2YVLOAmrTtXQSuoUa4FExtwO+JGYRX
SzrSC7Ddhc8LLDkES1ryNrEFn8DXLW9G0jaD3KXmleYo3rWMi3ewTv4VSbLaFnFMFailr7MUOnEe
vJJW9UTWldKxBKpD3+GN3j25cwkUPo+VLPCnjepkoE7AGUqZZM1H9qbpKisolinzgoGxwWOXw825
fhLQafWtNZwPesUXbGi0t9KUEn56X8go9Yu0l1G+3FPVe9vbDQ2JwpzKCtWtwuYJCD+u/6btbZWU
0jX3XMmuErIHRPOWHfCQ2kAj8tcoH+pVKm1wOPFL7QkDPdehYH0WbOmRE8fl/uEkw3WoUcnapdx3
J8lzrO/GnzZ1S/yzYXaPvL978KiImMkGLVeq3lIbI/AGt05tkbrrCky5yjwbmLqHI2KYbm0+pUFr
U3BkkXcHcdoVn5KmDmzKhp6Z1NMj0f5Z5Tkd0JhUp0USLDs8B0zpRZcfpL8CaCfOy4pScdhhmL7U
aYHBOgBmDLtk9QeZj2KwgXMQGmTZgGOVdROrbgoVBBrWYPqRNCatzMANuZyVeLyqLRupQ0d6LYZw
khHc1P8hHUX0YJh9OluiBu+CLQAcIdK1stVJfFwlNZG2ILl9udyY5ek/sFKYuCiiYkvLoFrGOe2e
dOIUMM9xszdNzrVgsGe93SoYDNFtN4iMi5NK8LpT0Tu8KBY2z0YAeakHDMW1ejNM/njRxzEwzs1C
lNQCcVYtwmyA6F1zivmtGq/XBu5YesejwoeSOe8B3++UTtN2dD3tQ8uXUcStiOKRKfMNYYZMKxo2
edJ6LWl4yYUC4J7YKcArKwuqy2Ds86tGYMGkUJCHPPFrbxGbVdYkCslCDwENgoinVzKvATRLJ981
1wc5+4drE4lSYSkWl6atMCBvtR8AQjChebDc0WGy7fXBT6tNbsitCDr7R4n9DOUL+j+b4boAu3Ze
jHcgcrwB4BrDEGk4mitRfsE5FTniuPQLagvMD710U5iCigNxyAUe04xeT2WMYLhARp0uGxDinvz+
iqCbPwDFghMz5tDGjvlyJgJaOrDGNxSrEdQu9SZDjpZ6X7vF6LhjnBFAcXsdZN93mZIFM30HoPFr
xImRVG1D4bsl/Pln4HTJWUeFEm4KbDPljn9HV6VefCBskUfCbdGa++MSBqVmFoujUikbZ/KcwUN+
7fs8yE9ovlj83GYPtnozYDjr6yZ7HzaMiKycLHAMhRby4gTxEVq97mG4iwQU3pk6ynljTYWN6RdH
8IRLV2PzhJq362bl/Al94qaEAwWuHWPWXpV+LV36PTBArQ55jrEbUl+jN7xNFCFJLluwAlwiKVq2
KysGmzG4j58szm+M81qHiCkeXNyROIAcILHlC0lQWLDUR2OqbowPDviL6TOY7F9uIh47GdKEobly
sx/CHtVcstRTd8EGUJ/gIGO39cgZFQJ7TqP/z+6FqNDl4is4Y3IQ0yaYwFCDFFn+H2PzqDBV1LgP
qxgaLQpe+qkESAvRxLIf46CLL13d64JiPAgi9KHuUVzCX2C+wGw7yT+ahH1CjoV6pURMyVn+MOoN
z0gZCQ9h0VC4rDeGsP8BijA/Yc+kPqQEGAO4qH8PlmLyPZO9MBAi2DaFklTGNkgoEWVXcOIM9L2v
YOfBeCE/wGqTZRAAukII8etbUl1y6qJU+oTTBxowDz7tDaEg4SNofGLFAXuGnf9g+QlSRpmAT/ri
FQa+HtD40rGf1d5ve6dKz7lw0CoI9LFQUwlRXuU1OJfIfmUtLaprpM3Zx9gWer303Cba97+Z5Dvz
KaApj412KhY0PCQWtiBNJLoPrTCI8Q8IDpuc0LhlbEYRshZ+coJ1Ev29p8ql3fiK4P623BBHTkLS
LAQdkJnzIpAftUvMLAITGf98GYyLIvyK71eRhchK8W3hDs6KEYbXDTp65yscYyHwSFITko41tt+0
8Oe15rTxuIsLHPBnhcXEl2oNoSFAL/HkHXVb0Me1bGb+oFjDxOjUVkV33wfEMfy3oHdz5JsAf4ub
LcpR3TvF5URiZbvgFVs8UDdLgLRa7ikeoqpxU3POqOAtrZmq+W6LuZxFuW60gEbyiPyiSULrcYZW
nIWxNF1+xi1+sOMYBu7T/qoa5iFrztC/bgx2mMTBIVXmoZ0KeMI2zCZ6Zsd5IPG2wafxvs0n5mdr
mLUwhFPS8c9UGmCFPRaRu9PS44wxoQ0SzdC1fArd9V83mxA9Yk7cp5O4HIo+W97f9G1DntqFE6pe
wHBZa3VgM7Cefn09ynauOD7S+BP5iY2DL1BNsuQ52a6nfYOb7P1O7GZZunXtMuc1cmFurjU8XJtZ
zdfQ/OS/fuIQeW8M5rWRsTcNpQ6kUHHwIUDv+VFEbWHnBx9UaQErRaP+0R+ytsm0Qu5XiT99NDGo
INciptTjQ9ES6D82AG+QIiazW5irLJtkNNVI5NedJ79eQjamrA2/5GzQOnoX+GQ5stcp2fvuGWHK
UaAqXmEAeG2no+ywJu6JC3Awsq4H/Jv4iGwVkoIDdGfdHJojOSqoH1ln4j5mGHim8H06UPwwhFf1
/p5Es1rJUy3Tr0IT9P0yZ2DqFuqhRj8UPrJVeBrcFj58yalCKo84cE3RqyK1vz7xVZNgceAbpcNJ
u5cuoCuJjbf6rsr99gmnMcJ/a2wXJDH2oDEThI+gDUL8bRg2mDsWnWJbjKAjZQ+Srb9FQ0BLcTyD
TPA+1s71BPAMuGYp7iylQnaQUj7CUUVV5uKBTDQHtPy9Cd81kJI7YaY9DmZc553C9Gp9uX8AJqNZ
RfWJZLPAdxu8K+6hFzcfQSFrf/ww0u9JdONsMtaEPxDEG+j4A44/46eshfl8Jr1u2syMermFzkEM
0HTJ17oMU9Giq+YCIYGM2CFxtzqqWL3im4XNzGUpGgCXrskbCMsCu3eUdiQRn7N6MpTfrIRfgZqh
NqHuAIFuZ/RmAfj5vm5u16rjDnaeqnb0ddOdVv5qVg+AxKptf4iUwM/kfDf6G/LRYyNEYmtvB5G3
ul+0e6CoSSpwsoiFN72YkaZaxTyQ2xTq2oJiioPYhim+6hpQnsdXeOXiqFL4hgqtUJqhxdrK08X9
PP70w7sUc1ofkz2wk5HVHy8iYS0BtSjVo8bzZjTwBdnPNCoY8/yaUUSvr7Z+L1Y+J06qi2jfvMTu
l52cjBOIQVEwxklkvrh8YIlTuno7M13wNGAu9iOtKgta23yu3QHYMRo85Hu2sPBikIsxbxsQh5G4
CldT0DEh+QNlPVPEzX3efNypkDNx+yJJJVN86F/q76N8uQZt442RazO1cQLFf0DWy8kfV8U9mcHl
Xybajcd+J2P88BgawHTi6j25HDGGwvkcK/1ny+eenyyMOZpz7bFkg49RlVMSLZE8UXT8CUqPW6hO
o/mrmjg1aRFoyCoj4ML7FFaNDZKJAToYtsEGt7Q2Rj1wtoTXlkE9WaR3GJ7ppgyDhFzpyyLT08F6
qh8AUVTARxkW0F1FjvFlRIClb83HSYNf1lnmNlG0slvY/KwoVW3mKi1mJQYcHRlpZKkNT96LLpKU
ZzbWDN8DKIpUarHnIU/TSxMwG4n1wB2V+xWyiMe/IShRAh7WxJTsNSKbe+qJpII0vhmAnUA2DKbb
ViKMTfkGkOLDOU0IvFaHLKs4hjOdWgVNLF0tb3SNALqSLxShXJ1CyZonNCzDmbn1B+v3sZDBsagp
+VS3vXzmtdPAgygBgg4PtF1vPYAfbxgvREBhbeOIZjP6BF7AmfWzLbEq+qqo460+Vt4MSCggOE4I
n3FEhcSNKa5o+3CipDIHWcl4a6t62G5ay9GmWZ+GrxfRRcVRIzZWWhbAMJDm0hoIN7ZQtliOVU4j
JEwtsbS03mve29yvMFEbp8MhK0VmbuothHQoblADEAPDhZUTgKHCq8MHfwAz8OWF9e585K6wYUP6
/xUXb1vJn+rVLiUXfd16n6XBHg/O5/QH+3LWostpLkXO4c++1oRG0btQFxraI6ojBBgRm/aM534c
DRIn35kHuT2p7uyDhgUInr/lJoFRykywwzoX+369/KxwWDgTQgoJ44BXDuhUG22RsJ5ZDA29ZM6M
/OtT4ekgxNGYuQxNWU5DIHvxfATLi9iSmgBjbt9eWtCNQkVtkQ5yCuZwgaGcogv1tjQ1takWaBYl
q7bcrtt9rvc2EBDxIhPtjFF+5MGjebwGFx/g5y4aOtfS+RMe08U06Tq4AdNaMNTW3MrLsSOhsDKg
7GeatpOzKjIPcZNco246yvxI1eW+7pAXzCZF+zMx/cIHhlBmtrpv3X8UCt32VEygRGASdQW8Kewm
yuFNJSrzAxXuCJP7v4VGxX7cNHpZgAIRmiPQUSX0uA0ozarMj16T549L+5UHTuLPSy1rhyWBUmA/
Dc2qayyQdxGzHGe7A+YRogjsCGjuKCgWROs/rnFo8TGrj9dJJpCv6IlglKDXv0SVLhYqnld5WpwO
+a9SbjaB7Apbv0/nHFhh7l2G4ddJWh7M2KcObjj0MwCLAh7RQ6L46sfjyAMKa6BAADV2LypcX2dQ
z58kysjeNnMbPE1DmvQrvNZf4VmZJemOGxgWUv/DXl9j9iULaHSqHXVRvUA2d7PC82QHUXBgHFFs
kB0cd5yUOH2aeVjTo3n7CL+1uSUmDQNJZpaebFoUtaVyHmsRTZIf+FUGjNqylyaRhi0sBCKF2yP4
JtM1b0pvau5H1tgyivQ39zTcL2YxLg7x/KQIT3lpH5XkQh8AOJDVfULpVJSsUIjA0YFaFdN9mWv5
XJuTHBGZv88KN2Rr3YjwYFmD1/7Kzmx9AQ62qbKbdXeLaJREmWqi0zkZsYjILCSup3roSweKHs21
7fTJ7VxdNAESdT7AuizOS4sKP2CA3fxTr6IA6XXdx8cCjq120GWALOZjDSzDqsAG5bWEpsuveU71
JBAqTlBz+xUPuiZaa1/45XWNBgtUxRTIDJFGkbB1Eu7Q8Ir+Ysumc0fHrPKXkQr77wVqQzMbs6sU
D+DfOJlhOG8QA7oXUTy7+UM/OB4q31l1qItpAsRgsbqsZ0oQUDdR7Ywxik8DTitb9FgGKQcwwOHq
6nucvPpOvk7DSQAytBeG7B9GZggc3eV665B7E9gnStRqJgKKsuzLInWw3wSYoU6pBoM5v4XXZORx
wq0oNR/PfsOplJ7uUmFZR9Af+oPsvUNyv8/onrede695bQyGPgYKStJrmX6TEZrJ77nP8FYiewxA
XhzF+T1hT1Fe5nddcFaHuUo/lEhOABLIsA139Qoy6ReVRv3viKxYe83iFBjsUN0SYtOzVk97sk15
TZdYqzidGxQ4SXtf0BG1v2SaSqXUt9tVwqk5sXcixMx5vLW6coeNA91x8aEK6upbB8XgVZV1VTo4
zZJfkkGjlgSw/lIKHQ+YRMPIY+cMDKOpQxAGExg2obN0cesaOsT/NbbT9xd5ObHRfo/vHcSMTK2X
7Ueo2CBR8rDKyjuOCzuiyYWLNZRaztX/U/gVsWBqoepK+s2fqkvSTsjcut477wTx+tyyilk4gt5O
9jhdYuCkMC4aN1DeRSncrewtdkQ5mCrynykSWev9YEaSChsu8UzxCtKu2ARyA/iz0ONrctwWRtBD
Mpl6k6hxQqP2RIR45aJ0nvg90dcp2sDkVwrE/4g7w9WoCbEY0qrFdiwSRorMehEGdycFjW8B3eGY
2NOa5/PczWcDeoU7KVhcAgYo6PqSmyLzJpCHphb4eCNmQ0W5/eW0ozWJWvh+SlxFlff/4xFy4q/t
UMlOy5yU+QO9kua+aMpGKLvXGkPa1A713sg234i1Z9CaRt1rwqvWr3CI8iWEolsOI5+ljYaEIKGX
So5oa8oJmzRjqF2//aOuXIKmxiboQn/YUwjJ1q5H5fyyzvGPRkaE0jO10ZXICr4zAjlyUmlUFv2k
KlQH/LjooB51oN6hSXaY6BZFc+rg9rnIyt7JT3SvKltPHzI9k6SBqZCbcoLbtajVfSdUlnpQ3KRm
6rt6EuxybnzsF6S5CNQi30Up7niEEB8qIB37f7YqUGo/kLALrmYRO0AQbVqXb3Nif4h1rQcOUdLv
cKh9277MH8YCGbHFPdmJC8V/otaXusP7Ch5T3Tl1bvgIW7bXKM2JzYIV1AZDOKd4ALcmXuxlJBvy
wJseulE+Eu0pwOy8WveC/C5xo5s9AP0BHJHorRHl752hFaPoXDrBGzhced7ISQWQhTS0qiACvdrn
mbu7nMU4RWkrW+gx1jOya8xZPNHrHxxyvtsJTtuf2S8khb+QAkjKiVwSwWFYyK1yXlcOS9QMoOwx
c6uTLyH+veXmr8ZJB3tH5waVLUV59/3ga6l/q4yeEMUbWtV2UFR2taKML01DQKt+ssVgdXql5EB3
BrSV0K8r5gymvpGAtpltgMtEmS8+FQctXo1q4pWrG5NYftCz4maSUDkAYbfkNpy/QcFpM1QEMx4Q
mZNGkVu0i0zHZ9NJJuFs+VEzjkhElG2qDhI5RUf6gSo2X3MWiMo/uqSN0q8RzmJTjls/xI8ke7rQ
cwIy5FLC905SUc4bIir7VkcMy8lMc6/ZYx6UbOFNVQXMV4IS3aiZfzij3vF6qEdB0GjF65oGzEC4
qplcMJadphqcUygJ/fpdhIN3e6sxQmjmXyf1wzDW7n/8B2+U9Q4n1J+8v+ytzwYVdEK+4fy+/Gn4
WTQNb9IdhHyNu6cHvCR2oAJ/skTksow+TOyPHLvHsgfbr0AfPAOTTVfjqDA0WOicmqrT4wE5PDDS
AptekDeUiagh9On5Dz0q6ZO+jyYC1hPYZw3lcNHjtXSFHBEl/COx5RGqm7PGeEteq06s699rgJE6
2uty8c6nAiPCDlo9apnP4p7clLGGtpP02RzysCaWbSVTkenkPaGwde6zWuArFxDqInSmk0lEcXpR
e/JTGZv2MAncLskRkIoYOG4oXzQcLHhGlS04gFlbKeD/ZzNKe1oF28poUG5XK7aUWXdPyK0OE5WE
SgzWIn2b42uHA6PQMGGqYYomt1JP8hizyoCEOFAZyXfCDupYg2aMD3Mc29u2eGJAC7FzaFFIey+Y
xnWZWpkWI2roNClsqKlf+Rh4COycKCpIR+eojFcA3cNDC9s5OCNFnIO+xZNbdix4Og5M2c4e9WQY
9ctGx/cC/x+f+PKXNLzf+7V03hrNQyKrIb0H0ETkZyH28Ye6py2Sn7Kb4hED43qFRwvOPR6E74Ys
imAuLW1uQnqWf0dgsfoGXasoRDBkTyUaBuYk8cz2udpMrP5wiQx2/ztReyrD/Swklq7wmLU+42WB
rQBdqez9jBEHOE0B2ztQygG8jUt67ntb2J/1WFCw7DW8GCS2dloVHtxNKsHXj6mLcNV7QggRpzsE
tFWSnKVTOR+989N9Vq+Tc1WeiubfFu1GgDj1sqZewtf5TPeYf1TfPVSfkyl9T+9cYL7Tq9pMD1M8
pLecDshFV4d60WEWVc6adM087gHfyI9qKmMmdUjk5KItsOpoBPJK41J6Sbo2DckUMN6sGizl+C6K
yWMDVMitli5aeOEsvKq9l7F6TyezGJB/g4Y8L15PDOgttwdzv7aSbgkIKVvS46lE/yo8rkL7GHmD
//tvYEzWE3+JU6yzsPSuKl0uOYwwrj5Hb7eSu53BxqPkndeq+EddnyZzzuVVFCpiTrE3xpKxdSQw
kc8GGZDHPMfiCiwBUe080DHO7+YiyXbjKHGtluwS+175ghoMLm65kbTeer44B1USs45+ggjU8DLA
1iQzWxu4OJZdAUYFNU8X625Ml48Iw90orNAuEV4FxUNaC1zvC99Dcv+OHxg3NK2rgKhuPGjKHup1
zhPr1+IY82XBbO3MJN8fPJXJ6RCIqHcyEtGAsp262DaeoObQY4Fh0MPRXWO05n6c0kQeTTaC6OYc
MhP7hoQhwkIj+TStRk8CLzuvwS3EF/+vZk+t5OwSjDfWixXaLGVmF08RuynyVTcTCQ9wWdbkrkzH
eB/XKQ+AwlzkdTuUzgfVrmXW8ZiAYjgbG8PjFw2HZTza94tisawDzsrqor62amzLnkJtmRCBQ5nu
xOpwx7tvGly9KLfOiKeNk7FOocGZVWjEvQEN/R6oxkRPvc7qjgMF5o1WP0x7l0uSDmtjqka2enVt
dPkki0tWXm0p2WdAmGy2EM6STmf6nUcI8XAkJ10J5mb9716HrmGAeeF6rsfWTQIF4HayNYA09iJa
VFaokFccfmcMJJYNqcMrnLlT2NoVm7DpJXFwB7LICPLChgh4/vXmrPwmFW86WkejFbyKn/HCclJF
uvM18MOrI3azb6lUAL/CC1Dof6XltsxSj8VyGbmXRuO4CKguxoYoWJePw/0pc8zi1dzP+c8DOpTN
zh2HFauOwGfjDFrr72OMXt/asdw3dN00VFxhrJUMm37ocfFpm2eRFJQjuvVSeg/jM64kQADGOMvZ
m/x5Ky3d3TjjgUqcfXEdAbso7Yh/CcFDkcO+h78MChiOOR1EWBXNpBbO/HorNzYL+QxfYB1hCiZ5
NnkgNxuNncbs5v4Li+Rue80Xmk4mALJOKGOkR0QkAZHHkdf9SOh4Ym3qO+1rOzDT5ADiwdC7mw3/
W9SSe9u87Y8+SBSvEbLi0fWANi9RjXgn5/A22CIyTj6UZLXdgezX90JmQ0CMZuEWw0mTLFLMU/5b
za3uaxgXhjBVDKowpRjn2yAImHgaZxgCGFyk32kZkEeG6Zp+97CbVXgyXhWcJ7j+YDsLcRly5FmD
T3j5EbDtnTJaJKKuzNxB9vM740otz9vAexGs/BpJbaT74erGBxTiGzUC2wQ8Yz0wCE7949rv6wvz
puyS+l3mTYMackG6R5cRitQNPQMQ8n0hrQELTK7UjPPV5+yTWufaSyP1EGEZUOwtJ8WZcu9CpQCN
cOvzcLMbDBuZrYv24cV+oj9quZ8ZLCAzB9nGCnZU/wjz09guTDhY3nWk6i3wMUaGXWaqWgcyB1HX
w01p8a3Yvg323m7E3YPOh/mh00Qrx0S0clyCk0fN4k1OdhlMCCdMfImIrwVbfNauFaJG2nMBC7Rw
490OGL4VqS9z4goec0YIOQ6HIwoOuHlYTh9/KspmIOkntGnagQT2BrCIolYNz5svmGOoaioDMvUu
/oIYI9h2RNXBMBjuVY3dWHqmwa72jhlFzKbzRda/HpZ6MccUk6BB7r5wrghD2yxRv4BOLV7xunvb
K2s7LwuZJ3hT9jzPpWbdITq81wRvyoXIXIIUtqXxY/LQ+b5IT9dniDJT/m4gREqsydzTHKq7rY9P
CivASu7fESz9ioMeX8PyeYsgfm5iXU5mknEnRQ7HjZVr6GfxhV80ld9vPp/Qsw2RUsSMULNyWsTH
VDl3cbeEpOIQblU93OVa6xUFN4D1boQDsKKaOkMGh/616Ij9Qt+e7OWQEz81YRsNh4hNFFKIaAXu
iAr2UmvdVkKKPYAs7AyOj3MUy2WD9ImyLYV/HgZ7NusoLcbs0ahemqt8QIzcY5c4CA3I9oxFNCA/
LMPxpU+TA9XnHbkvgzIOUvsUbrctiRq2g+6MtgVQJaMYzu0kJkEy03/5hub4snulAXGwZYHUcgf6
ogv19n6tHezBSXmprEBQBX8flfReD7OMjplT/d90ILx7Sk/YmA4xKE4jNMt2zgd7//mD/u1xPPEs
+SypfUmGmOM4FOdHvAHNWmKmqGTpzIqIJOFSXKFVvpJtNihg2Ynjk9FJrtUFAXfQHbFlcBJtYmbn
okYgCHUcwRegz1mWmbG0KRY+Df2sHXRgAAD2+y3J30FYQh1/Gjr0e+g6gJav7eJEzAXE6Mg5EgOE
NB0f4gs+0PFoS3TnJ0yQCinn2G5S1tWQrYlI0ydTMknAbmRaMWVFqhMhZnJ1wPt+LUT80eNfvwbH
1z3eWqZ+Dba/BdMlU9Il1E7puwRYPoj1T8uK8qeNJ0sMSlcF/QWq8YlQhL49hY5QtKpDtuLEb8AW
EvGVZdYoFS6TVRwNsskdPwtoEtyXPjQJED2c5UA3W6mr4J3kbnPW4pFTZeHJsN0AIG//gFFEFvmM
r6WLctxiqx/OFIHyufzK3A6bY41V1NhCsaytfIHElSGHEWAH29e4YouVwV6TAJ2eGs2dL5scrITv
/gDpYH9yfC4A3+CyiWcHBXcTxmoo44Qcr6+yG36DV5fzH9GUmPBqq96vqjCYLahxSDhxZIk6xqf/
+Dx7iQugjZXFddlJnnBgpzmgKctCMHUWaFuLyqbvSCwPSR+JhQNBqLITtR8qOWm4jAUSthji253/
bwUJhLk17RbtXtd2aR3BEFXy6c1HghPL5+N/4fuVQ3FzP1b6QpG7E/XnC+85qhUfkI3ucAzbmrQF
0pfy3QO6V0Tys2jlUcj4nwRXq19l7B1twX+UjryuBYrgKUpxhPrNg6aMVDzZ3mWiTt4knbNZ3wzK
tAb3gQCoYiMrJ5ZSNZLUsvRyGND3D8Bt7AYcnIUZNKpYeyndqK8sj/Ova3gGNwt0isFgdyv+kaw3
zwd44mSWh0W+SmBgmze2PmAreSAsU1O1rznnGd67sRI8OxwkBRmWyJYDdE5zEhgfov5AK/fBmmWL
alGnIadC0of3g4koAIZGgdrtH58OHDBaXCqghtpR+qMLEx61NDLx3kvH86DHEPi5L5n8Q5LGto9k
cLVEhzeeFQRqIeVE+XcCnDas2P+F+NfnruWS40+5GluVgDgXfDIsc9B71StpUOe/AFd+CJTYqy9B
bv/H1CwEGIJBkLNjelPj6JSkGdXSeoGylxXGcoFUVzBiIth07DSdzHQzhb2ZuVX4WfAB9/46OtVj
x6YraHC7iZggyNs7i8pABBPcq6D7e1TEYd9xAYfS63Qyx3BLPOHir6gge/D4fgvSxZJRA2kSw630
XYWg+MxCmjSdyV8FLy7P6HBtT8zWssVGI950s39/KOTfQIJtZ06S0JnjMJQXK/XqsbBqD+uEa9dN
hlHpLi9RVKW899V3p9+q5FqoOFVrEJGLfzmbIqOLGDSY/2oAct9tykTm9zmBHSCOFbr0Rv3+66gF
1qohkFzdVJHp1exLJ2JrhvHBaQgHn1c+JoZ6hZt9G0SMduxbOQ4pz//1N3j9RQ2FjUf2woJaKdtx
v7r/yB+JzOdnBR0ty0hzVDn/G84Lr1UzWmZs6bpIdE+AVqfY1gzicQYhiog8ly0QpLfgbOXh+X70
xf2+EB6TmePi/DSd6Rg3SZq/y0RQ1tbWdJUNxIES4Gcd61tgYzl/WV+qyrLC8FdmDd0zN8bEvxrq
bF6cpkQ3XFQf0OTyFF1mqjuBfaHWoKGmX/zWYIsE2swmPkIfe6YQOf3Bg378mQb2qtx/4uIIvKDF
NdDqD0h418y17zDN/HQ41+Kqe6q5TGRWLlCteTGSK8qbTWuRmbqfT1Y1aCnWgjeeplh+aak8vP9q
fdmtjHwOps+Z+XU4scDoFtla+TwBez6PcN6dM1YZNPODOoJG5Arjc+EoJCwd3RqmdEX+bkFbSwRe
spw7Q4FQCwB7NSF1cG8mkTA1sv+GWMjVAtePYTZHmBX55KmDImALpLiZchp1CYEIJs4ml3P6mnk2
c6TI0ipUFhB+l4HJALuqc/CT7nVZL5bc5QjBTjWRwm/DTkHU2gqwDhX6sB2lIs4u/789uVFEpG4m
HjE2hU3SWt+fwD2Q66eTOL1ourdrIjSDpVooKJgXS2fWH+M3JU5t7QSsuzILGGzJoPwJ3GVi2k/x
deu1ruDfg3/RZ5eLjUAjAORAaUPQW0Ghu3QwZWVuNxm0ML6C+9QhLHDu7tK66W6bddkkTMPWQBlm
5KcQU1zVc2ElCBYGlCbCBbUKIXEKhOijjE+hA8edL9hEyRGto6CKpyo7OQZ4EcOw3Vz2XesXcEBL
pB/hmvcoTVQIJxzcMIED0I5piFVtHReMVWJyCkM1RkaejkQTox2W5UY/jU7IZefjwvxqN2jdeejb
Fz0/rdACfhpbEoVBSFsWboRU4GWfgeva4vgS5AFBoLpEu3+Tu10/IsbjumRmf6N1bnN5XID0+3jF
faXPN2OKI9LiLzLmDIHAYk1gpa6a27Jt9mcTQf+1oB2G4kO9AyWybPveE+JbuyPYvbH+SHg1Bgc6
4Je/7h2d8ykmN4WlB9+3YahpiWdrnM4KFcOLaN7f/I1ZvW/bJ2m5tmEDA7rQSQdChhEp0gcW6qb8
rl5P5gQOf1oWGSObMbezdn+Xtw6FgiCCAVRJkhKqKy+7pVG4ImTflKeLtj3mkms/jXWDFXQpTUlL
5wI50nMJGJ9UoQQXZK2mL3PhY4igTUNE44Rg2RMWgz84QABvibqRV4nOw7KPwsU88vsy1qZVhZJf
Apg5y1xjLGl8dTvbR88F6rBXEWf4qcjR1aiAOe8lsLs76X/WSGyRj3E/zgLxMVxwwe6kMwNP9T7K
Zep/SBppnobjMbOCaHVAbKGIiur3X7rw+RNBXMEgQaoeyrMJb9vnG3BCONOMPxS9G18FQGlefdjC
uvmVc0QHrJfRSADa8IZeR2m/l2NSqz/w0D/k6mN3hNzsI/KSzOo6GhRPKiQpnXjEBsPqWyNmskMF
L3ZQoY0uiI0QRTyF9Ef5VOHV4ZYCxyRZOplQPWq6rHy21TRbvgz0D9dM8VT/rRhyvUlGqvofIl7N
TTXuWf5weDRwdGbO953Hzu75LbLGTG14+8LIb9UGdm4KXWnDyS19acZ1qEDT0DpcEertWQbkdym4
X57GfMQYkEcP2Q4wlcgJKIp4j9i2kpdQA/B5z7zWP4D5pti7dkYmFonz+ypZRi7EpsXMFa2Hae2l
c+s9Kr1uwJLJtbyBEZHvl83lxcsSnT/p7OTngCAzVp5UPWoLmM1RHrfvy1sK0/bvwsF8xKypjN4T
oevRN1Ad9ztQLfskHup4cir9olG2UMvFDb3pSamH4sJai9/Iw0WqJbdovNtLpvawnnPX5DFREwaa
Cnfl2KpDR1CriilNEtew5VeLQg/bjB52TUrMipBYk/pRbNbCjZEyayhUUxH48KoH2WEYw5TirD2y
t6Jz0J7b4NdtFFlz7I/J0UmL58R/7OsEYdId4fAWc1bVfsZaMZwz1aVdCjtoyRbVzQ5lEw3jh/P1
8GOBycR4lfUAHRtyR3yIOEymeq5bNDXul54bfBIi4srAOR26iATF07TeSz2K5ma9+WmM2dj20sil
3Xfigl26BXuiEQHM4IewwkH8QixOJgUYAcNUqi/VJMb6e2IKzjGR+4L2zePNBZlyk7G732Sg3tFF
9UE5hMX40W99a7S4eaRf47EI2XbxzFveyLwJdIVv4rSiIVf7z+IsIrpszXU49VPNv0aM1od+M2oY
M5MguXM2JdtQCTevIm/nPUPB8GMUgqWmkVMR3dg2C7CwjWOoiGKZ+vFcXywdo5WjB9nVtwA5EQJe
XQbOP50V9TJrLamgNuqpM2C/8AK67VhuflURYZ2H8G4tBf0ZdTF6ntxVTygFXLyn96pNhCkevgfG
qBjIemFT4x5ZT/i3YBoflvVkSRwvvf2RW89UFTaNNXH2G8rYVRg3kLlWivnuPwUmwKPww4Fb+Ha0
7PZfiY6HjUZ2JIWuyPGYlS19iSRUQplku1L/yMZbLw8UyQZKuRoODGGce/TC0VeCwztyEvbviSd4
QDszFGDmWTHqMBxKshyIIyLRUZ+xtnegT+ADSGqaA90dkxpizi/Je9er6mvCyHg2mFQMKiGb3F2C
8yc2I/W74/hKEh98D9heA5MpLN/ujzSEhJqrLFfafoBTGrxYRBL6FHuymMxlt4ojKbt1lYlaQSJs
70thYkekd2MNnzdF4iz8JA4CqY4pq1WX3dCxalZ2bzFjVh2xHOLlb55jYmY6MprHAT3FBAJp+DLu
/ufCsXishAWcYHlpR2e7vQTCmGjyixgcPitY6TIY0J5hI4UdEdOMzjIYqNIDcATGKzEpseyYqNHc
s0QNjce3YY53UM2qjW6/qRn9QMtA1BXZM0Z5GGuysr1XoaH9j+OSUcgZhdl+QfmZp/qhQApUVZ6N
UITB7/6PzsW8YvhVFe6GXBC2KOcLpRv5TUKxnEzClQB9sUJEnpg0n5JvCKIkjW7HhTrIUlLzOpiU
dXw4UFJfKQsT5Aj5Mnku6TRM2BPGOrfCvQH0ynwoRXnYYvbfD208E1B9Sx318AbfFryjL1J9Tbcw
QSc1z57/tV5E3LnucMBEiStNxG9TGa7xqcn+vrlt+SvpSZcHYNGIhH4VwRQT2cYcjRSfCCSSp0Pr
iWXM4i7bnLh9KS50drSL6oHnC7bnoFdcc/ld/ADMngUzlMproVmE6/Wi8bsFZ9U/uqcM5SlgnvGB
61yOxIUeEYBKhdUv3FnJFv4HkG6k0AC62XgcRbqhueAKbSufqHEgBwFltnY3Rf4R52qgMJ1YmosF
MZZvE0VzYc4KVTNOVAGBfubBaAwxgVvgzxWPC9ruQO4+ExUMUtkFKQGu4a2d3EcENhgBdmDSlbfq
J4YwZ/jczYjDbjYZoqL69CCOvwjDgOzbxUPPlo2Nn40sQG3fU+6VWgONzTUevYQd8Q5Kqg0rdnYR
7afptuQ8rcVDMcM0Bkj0PRSBuPQHFBq/TPdi3lsudwm55Wo/xt3IqWWXemTiLDty5mC8K/H805h2
3vrF47Zt+y4oazzLAw5mlN6qxQ52Ioz3lk2arquTTWkNKzFnGJuon0U1/0avwQBooScw/T5EXE8S
h2nfueFwbfHBzKPi/JAr5piu9+OAcbWhaTwPlcbWE4Mj8IRKkqfKuZqFemXZPzv0XaA5Ii4obKK/
b2uWMrrmOta2JzVcRsPeUoGMtpwI+YlzlDskZmy4eTI+S9Yfp9KexlfrWw5yDTFiz0Xs62hHCRrg
Ua8bRQiHC30rPz5vH0Ml79Ir2ooxP3JtjT3056qMmAfEZ3m5BANNHbYtZu1Xmyg5NQdmjAuSwrkP
bgvm5gOdZ18w4quBfLXWXQwi9AlPxlt1I6pBzytRvK7h7OyYzUdxvYaWwgUigYs/jgMVX4LmNZHH
HaaGi9+fukIReVJ7jBKOcHf8gGCTQVHTbkWrw6vMtOFt1Fj9gcWJFw9tDznUHRsyQLhekV+UZyT1
BZwsFEUXlgnHGNrvkgdAH2CKsPHLGjdxMxvrUMw2refOLxNhfEHKTaLz0Epv6Pd3UF1zT8rOMJeL
GBobaXOk03/jtE1bDtH99xIvySNyYnY/2xKpAm9zb+pCrvOEY79i5PPjf3qg9FtlOpil4YI+U2nT
2D0wJYvIX7eTyNmjLr/vSQV0gJ0/RwFzoxbpgSJ+hNrs6kP1tJOmMF6uYKcMbfxiVD1lkLNVoo8j
yV/lgxGiA+B+sxO1gHfWyPv4ar5IR0O3H/iGm3QPdimiLsOirKE8RqbqoKyfASMfJ49/J1UqAHCn
SCiamlI8V/iAzzfuoqnEmrHwMsh0WW7kTaMwemc5ltH6Pfr5FqiyrW2Hxp/ksituUgzyLUMAO8SI
8HJ/c9jYj4rzBXPzvZh+3qNVnvBqy0q8wh9kFPK+K77NXMAuAIpqW9TOvNC9WUgthc+ZYmmdQMX3
wKdbMOqTGpIiJlJLuA0S1hjbGnkMUxsO+hFjJEO4aQajXxYWFgdcRvEWF8k/4iBOvqyHnciT2xVk
IyhT2JNZf6G9SWzpbteSQvNNJXkytBr+DX6+8zpYfZhSThzD8b1CHy+LB/nB8CnvP1/GQipwdCcs
McwZWg8i4lTM9OD8fd0uPW5VwHZ9B2AYc8Q8xOf4Entik1WobUqUfNGkB2PO6zLKX3coXUTPBvl0
k17EzTzPD7rnRu8MKtocxkHEs0xh/AldL4YsSvSM9/JXOS3LFV9Yi+jGDdkFZw0YJg53IdHpdWGo
SSQ+vRlKjCPEup0Iq2VfCzL2l6BSDqeqm7EzCX/KArG4XNQDodCeuqt7SlduPxRd6VqJ7ugfR1ve
iB07Q4XBMom++YF9IFEhgFvWnf2025Coau8Rx830LuToicDZxO75OJl5sc+Z+QAjgjMLTQaxwSHS
x6gu+DfCHaY5CrPxNLjFTee1Wj7aYf/ntSfPyFZ2fyDwYvZLBTZ2GO2ekwVb9aO5qKfVzGj1QrcU
DkTmR6PH0NfMCtjAEmcFD8Her2STxK1g6dR2ofAJQf/Px291P60ViuucuGvuzUtwXhD5iUknsGgI
tt6bUSjCm1Z757Cnlvqml+06oamRjJRL2lPV5yAWs/saCcW0GyNJbiw71TdmKbA4pSO6bNPf3I8R
QmZdmuacC7kMNbUJyokbEJmjWWHLhc7CPfDpIFlepVYU/GaY63COdRevTISDfDZSpXCLqAuHxBBo
7vS7XVlkHkRBdeaux5Ji0Z5Hp5BqK121TlJiFztZoA64tdsqlF9XsemTtYbGGJk8320VrVv7+D+K
ZxWMMs3gTzRDntt177SgNVg9mrwddK1wmC8ez2XAO8/dvfx92PVY3pUTN8l0PmXlYbjzg87Q3Q3C
UR0mI1wQO5zcjQ6KkNZJObLxLdIrDsZ6f75xJOO75kU7669yldD/jKFewucbT9hMvv25iNvSua6K
uQd786DhViCVtvRdt9ifowjdDvJCC72RdhPyQf6mw9+dLaP12rKVKVL8cN2Rw4SuggdUA3C9a727
DR/6zLLR+JcdhAooTdLnagpwoDMXgkSqNnxpyC4XCWYAbsskPvRTap22cawTfNRlY7JHp7389z/G
KT5/jP251ysHGCqXHvLwS1TcL7oYz+T9iSNJ4l2OJhuLw0HSimHxhWvGGZSCQQq7oUvDF/9CAsBL
4k7SZsOwxGE1s4JaSAnq0Wji1yBer+a2ka5Fy0bCUeVTMmg9NG6Kmohli8DUA5yow/HsgcJ+hsWJ
Uz2vAbHRW2YhmMmuHRXsG/kCoMv5TDdtlDcmOY/vr1L+lQjdBe+1viCnSv8X6y3znZx20C41hfzA
ryyipuODtZbU5fVbzJXgR7kKpQ+9Nlsi47vNOWZj5JL5HFkMqa/l2YmH5vf8kXBj9NQpK4Zcsbdc
bMMgvLVaKUFqRxF7fHFTNjK5s7zduPVbVLPE48ayE4rqXNSN5Vzwx9UZrQ5z+otrRTxEgC4/JnW2
GzC0f+xoXvgvJcI7hpeM/Oo0GMPtwvgUqZ7knzNcimNP6CSPggybRk0VIvMf5j8n5Z1rlLAIPf5r
AVRAK2t4efhvKmke10OVqK7XqnNDmAyDq9c3U8RSBxcpombZL5ABmjlmtiLpjIQZC+FBX8mlM2Yo
SJ4mgeJ+R+KW1DRiTqxU9gW6tf18rp7XHyZuzhIsjDhj+VQfTw4YIo5FYgluHCQr3QmDz13GHpFS
AVVKD96J34YpSU3thiTt9kLdqcio/8oMWxC2nzKawlwA/k/7djLcQLW8cQtbkJOfBfvJ8984DQfL
sBL/aZUSRFHYX5HyMD1ksLdOXbqzHgTZmz0rlsRVlqIQ+ryVN5vBH3WbE30UURJZ3XBFIfy+X9Cg
4x/IRhEEhAkI8idWDHoHxRrv+2zfULWmpCSt68KtUrSwTgjwr84d8ndzsHwnkDijD9xCOy5+Sz8Z
cbf15/fanwq9W6O0LPLtVj2Q7YDCQmqXOAT8pj3OuQF7KA/MzghQgZA9dVqzIgEg9V/WClevK3s4
EZp/8a4PBSwLolnVm0fEEaCJdkUEeriV4XPE0Bj6/eEe0YnQj64RCK6pXhdigEpNOdDEGfHjC4e+
0Lpg9FlyyQCLc2CdaSWaOFNqlCGCwcMX0NIYXvl9+6u7HWt05e4r2/SZZ1cROXQOmLlyNrROkKg1
z838WGtvsGLLbZD9HlljG5J/ofrNyL0GjcWvFzpsCCgk7wt0/zBtvJFcAiT3hFAPEnVh6dT/Kf5K
n0JpEJ9zdX90c89Pd7ESTf6RSocsfmjnPhMba1RlsVRyT5AzspcbPIHRBtvlz2sq62FnjPdMJdtn
2laLojTp7W4u2/eFlop3Pso7/7oce0bcAqps0Q+yz/A3FqfndMG/w4CjCaPl+ik8822drRoioj5+
FmFtZc/823sfUUg61tbBGTezi/SjDqNxc1OvCZAJSaQA7JwOPsQExJckXeOWdpIWhEg0tN9EwhNU
QT80EBr0U9jjVwxLSXoxfLm/FEBp0LTIDucfNkHETm5WVUdV9SJ5q4sQ42AY+Z6r2Wq8bxGj2wMy
+OjPvgiMsGW/wXAAaSPkvFmT2pow9qwGX9n50HVVeM2PerpUXIVxCofknlqQYkzqbD2lzy9046xT
+nOYrbzpB/aPW2NXEHZwzvS9RjF+JMA9s3yIF6+UVEGrfUzGhNL+enk9IqXqxZYtaxK3j6V494Eq
eJcqCD6MClyum07jEdWBP6ofXUbMfRQr+N748T5XbFRcHk07AegJ6gBoC0l5kwdmFicKpGbiTqWP
8ElK9Z5RZPzPYd01AVFTtsosLFlj5nlrqa22HQ2v9Xjw5j1/bSXHbMRGHxONnowUEXoCyV/E9TFB
Lgd5VriCspo+BUVyA93LVl1imCMj1Ry/ot3zbfWAo+1mXF6kDZWbP/DWj6A/MzB6sVgsvOgNiOyu
Fx0NnXd0mhnael5L7EconcyN3ch4vtDzo/jFJWGaz3n/IgIMna6BgZ/hRndg8bE/PPVb45+jV+vY
xz9VDn3ek5TtJf0RwJEHkk/tV5/qfi789fQ8YZpwydgfZxJwu05g3UwqTCw/MbNBoVrik1j8vFqz
Nhh915lLazYPreXfmpVfiAFbd2dlcWHCe0GUREl+mbtubLvZMTvsePmBVe0kVWYoaup1Tdb/SnaS
DRVWO4xCQ+2sz2mQ9wcw2VNp6Hzyz76HXVqClUu7Q8IPndSzItO73V2ysUVnn2j08ZHGncXRAI4H
2Z6fQoldS6R7mEyT/+ur6cr0Aw1IfyvztmJN6LG8BQC+IweITI7U+ZkwzIgQ4flSTCVelOk4YvsG
b3pB7J0EPO4AxT8Y0Jb2o9/gqx35ZqoTZxCBkbwPNPsJJW7CIZsOZ1eisXrsySXAVQ2DEthx7ZZ2
rJc582IDfsYi9QI7DDxVWW5bPbOF/8xNq3COf9VcyVdSzTy3NYzgPSagS6y+3IkLnHNmYVpQG1Mv
FfQ/BkzrK87/9oVjBUJJYiHmK32eKKxwwJDu9GndHhOH/Gxf9xl3tMaE+mBl17xJ4vvAeuipbbz3
ojw1xR8Z4UdkXnnkr2h/SLAyCZ8+5WjPoZhxXtBC7lBR7E7pUBICedph4ASLZHgjQYEinnF+2uB4
/p/zKw2UlgtQVPg2i+eCeFyRxu5k+xPpFmPEKkj6mDDczjK1zs0JKoaCdCbIsHBpeQ7CYX1nXuaQ
posOg+EtlPunanzC7DR449NsNOkXFQXA0vu90f1bYgs62cu3E0FpXOk1DWDOici4B9RMamhTRqvM
3nOlcACFeQJucLx3tv9MKEmgWQzOBurgDzIyTwlTuAYgnMjW9yNZ+JgmUd61QW/sYY9RYlxvOYbA
4685eDQ3RVanXitd8mQ6nINu0HAXGE+r2dnwiFjEZQIwwzRjMz6aGPo8fXDKRe/x7LJXcKGYtZhf
3pq9aKsqrNwmHDhpHUFaK4n+Ew/8jTnf3v2CJItNGSiliKnPObjeruvLD4GhU3rX8DZNKcKhJzd6
7rsZt2NePvm0kKYa0CKWB12MR36upN78MgLRcaH8B/aNLizkFFDKre1Y8HeycOKkgrxh2xUBMht7
M2tbZvZv6gIsLaw88qbr87/wx9FNth90NRXM/BBXaw8e5dVWXkFyWtwPgzqt0Lk+8GegDY626uof
QLL5EPzZt9HSLvSGSvXpClH3ulND7VUS/mAkmnn9Q8cCFMRhKUsj0wrKMTJPSGiX5auCFPaebvSv
zU8Ov4ZaSSim5/C2bIG5/j0Sw+NOzQzHl4YB8F/ytlKFWLQ3UoQ4jZBSrKBV7v4AGJpwoaEKrqtf
h7AhIH9S+vORmq+uLnDV6UaBFUCzHPn/4JsPOQLLsYI2BVPwyO2g2RMwNv9Ff4qpi/zEjoUUBbOJ
08+haTdfmA82bsO2fV7EwTuO1QGPCxqlPZaSU8l+R+jViTlxrZ+shf6syjUGQHofmVu7M7FTSJAp
2ZI4RhD/k8auEMdGdIgFN43Lp247+2b9OC52IGo1iCg1BPKCTO85+Qxz3h3ZS7hVfPZ40zRDdcC9
JIbJazEPPkDj0kqGCvWXyOg1fGJxhFAQ0yT+bkwtLNNYEbxGaYyTa83lP6qNePgOBBzwxZYHu2mb
0LcJqPPKto/+hvifkax9EBrBhIaUkoFPRBkMTin0y1abgrfM7bOJigAmdkJO9i30kOridSw8EtxT
UDkhPKjurFqRurNYZv2mhexB/8kGIfQz0WkOge/PFNe90k6sSlx0XxvAJIHxBpi17D7J+dypV1oK
bgXFE7rHtPVaeGhCsfXxQxSANtq4sVjakJSv2J0ayymQXDOediQryT2YWXqePRWaity/1y7FkOJ6
T/EeOmv83q7QsqHRtWhr2RMhxeiI3+3J+CrwLRa3qrUkEjGlP1Wimc8i1CKA3zcRdKxKCnOXYC1s
u+lf7FSC1xuQu9yz+qyt5OH1yAnI45GPKnlHx/tEVAuo1Quu6iz3F4Ph82NyL/QuBpDq2R/WCbgc
TxpjDlRTVy6x5N4wsO67OXmFTsDcPICuXgvJ8VRNiZj+Hd4e/aa/gSxK0v+PA3IiKoTwVPsPgHJ3
I7JAiFLnh/IZgiMgRZXRNWRm6toBMRqzuGX8PqV3zJ/SYn83rgejTGPAcvwwq836YCr7EZpFFwr4
XN4kOzLrFK84rFZfkopBwj9c/Uzs+Ro/oTX8UuD7fh1aH9kfzc0UKr26vIedcnW3AXQS/3/IB5Gy
SbbAwWEnMTA+UWGH3kWZ/RG/t0rC9VcBomsMG+gfidCIvDfQi0QlfZ+sMaLfN4/sXvUZFiu9coJL
QMA2UzaHQJDKF7B4GqrkCTHNDMgJuwjJbMb91RCSx1jByVaanYQr/61FXHuwgidPZsr4d8oCkieX
xM1a03uAKPBb97u7TGRq4Vt3On8FFsI/R32LcBfRA+ACr2BpgHT7laWnPo6whMdRZ0Tsn8OwpSLB
S/WslSKlz3ZspEizY5oMkhfKb90KwbGLMJNG2002bf2wYcOeNf3HX5QZdDoC7pghgRpWFEjkR8MV
vI5Jvgw1ttgbw7YvvTydOb/d48DvBPGAOGzYPK9/15UDmFmyAXMr96hzX82r+0C1yNcttU5FvD5c
UV9wR41gPQst4+N+zIA3w9OUFLj4ARz1+JlJp2P4Wo6fpqF4LeMWHYOTMF7U4zevSBI+HqctqHKd
746vNG0PV3GXg0JPOsOHmDslii1HhCzELRadQ7TNx6zqM8nV3a9Bbxey3WxaDoC72OkfD6WFsSfj
z4UcZjkHaRvzK/WLD5dsJEN3qGeii/NMMJEAQFW1k3uwki8SBRYRL+V5VbK1AHZV3ags4KsSbQjK
n5gq+4L2BkHj5ZEt63f+XKdV+97J5jfxQxhxnLjXxALZPT2WESOerWT8FacoD0zbsN2L2e0aCSXM
Dsi7WRvlxYlVwNryu1ZqfrCxeiqUQ9CI0cRYcIchZUfHTP/f+TEP4FnO8EzeoQtLkrKHPm32WgxP
V+xgNXr/ZOzgrB/b2ePqR2B0CGfzfehkmOxo8Q0pr8rCdwYDbGMR+BonH/ImpQAwkxsIcCNATLrO
4wCnOxgMV1iG1zJTWF5vC3gFyHY2G9EW4zF1UEPrhJqaXBeV9EGieF9q1aIflxtnNVeJK0ytgNc4
JH/FuRvEi0bH8T/y2xMtE2SQZLoegBAkBhaFRaSOKrf07S9lgUSyHeltNBLLXUMAsPtXrOk2UplK
Sz2V32DQcF6pXRuuztZ1jtPjUjXvLKCGWNA0WTzUfyf9UgfICXoyz0u8CrtWq4YPN68tbV8/705x
aq4YILh/pGDKya63mEyAZH6jsi6VLUmYnoqWwt9gEx/v2OynKd+o8b5Z5jfrBgKzqqpG7VvxovVq
Ihwa3I/hLFr1vZsJX/TNfH6Y2elYDQfeCCDB/V5h0/96/X2aGf8TuzeLRqv+6Py/PY4kfaIwBpvz
keWLHCC/gi8jmxvST9AahfpLUntKmFr43p1Lbf7PWdXGfHcLrfUnJhExmWQq1NMLZ3asPiUdimpa
0j+OhXAnUi/8eEw8+d9wPEG9u0C5mqQbmpFTQ0BZebi7rEBLNhrKu8XmWXWCzy8KE20bg32Ss65f
JDtFGN1LU8X7tzR4Go4187EVvTmCFkqFi+nrK6UizsIk2/xwZfhkrL0yRpSaKDA++tbKl+BxLVvQ
k88CsKWf8dn+YwhLUMRK+Y0PHgG1qiFW5cc+r5sLkMFoJNPhXyk3xC6A2CJK5ZmGEARf3WWTtZQ/
ZF5mpJrdhOtisqCjRZDoPXB9KF8Rq4F5PdnrQ8UbhfCzr0kDCGpa2kmEjjaJTyyQJqru81Myb4v8
cW7DZO0Gx7kbxfrUAL96TaoJXXpnY2jJ4m1p3DIhs6xW+w0uiAJvWslgPYbfZPrqGpMXtU0YQKgA
5W0BIzZzvLL9QYR1yqpISHhLXso8Dx2rYiadOknsmXUNAGPAQPiLKvopOFE1AA5EmXGKv7zNNCzT
FBD08eMtRdthUFVE1kL/OW0/Asifg/qmVjWyaA/ghcyM4tJOQNC/X7RiDwoe34TPWE7HDkbf6alS
UuqlYJ1OlRSgPZklfVyiP49GXK3WLRhPeaMmWqDmkilYtuR4S3Pda10R3zTgBEkC9KVZ7cBTRZyo
GpAyNotZgzLOEPdGpIeOd2ZxMPQEPiZ+4jOi850omqDDgxwr8GP3Ju8/fcnZ43joig8ZKbr1W2SI
uJJKbJoVXbqJ0KMIO/zygmjdKtYI2qF3wXw0aZCS18O0CNklnYj4RNb9aG/1aJQAD39RewTvUB0Q
HErrQH1Nsq51zEJ+i6qNQNVPH/KQjKbsAR/Ad7jOPUmivC+IMzimkviCYKxnlL8ZsOyA1n/J3fQf
tm9aF1UUH45tBkCTzj5cIvNe6oj9Uiff5ITrTqVTqhEea+C5x3fnjf/Far20nmaWYU5Db05Ktvkq
K/Ddehl+x2XifPchWq6SdERYFBNFlepeMEWJrBjdHgbFTGYE1S6KI4GquvfT/5/qjQ2SylETpD5b
icixPsw624IrCQxthcQ9mBR8lWORiKrmDlsxwDgsrW3O1/qZBGOxXHbIpIabyJeRS6PGBBtZzWmE
VrW7ca7kA2btAcIZQAaFEmfzS+XacChs3EfGOfncoef1YbJkvNAPf+bT9xn4JzEf4Vdd3mm1z/uW
egn/e+qT60syovoJyPtNzswxoGsXvOah6ihYMciaQ3JtQ7hwwluRZ6dzeOtrSCXUDkHnvc29mttm
+7e6qcqCSE95DWUZCxezGZqH3y0BX1AGQbt+/GPOyUv3j14yhiGfogj8d+4Eu51OYOyaEWh/7aoz
4KtIUcUd1vLKqK/Qh15vjJNxLJBFDxnBU7sdaHYALhjajbxz6UBVO2w4pmOXShpSBmuMfwqNDPOX
NaTEkHeKGfVe/wYOB7hEunNF9wZXaz69eUnK9uM4kAJdGrIktAIGuBIYm6RUOm0OU0p1dlsJMhGb
LrOt4DnLp72ZrFNInsAgEbq5Tc+F8pTaGRchur1I3bBsQB8jUnDdPqTmtbcig8oqRTd6YutjjRsY
YVzTvz/+hPEOZD15uSoWIe1A1cLXuJxlJqkSm1d390MBSyPG8pxDBslGBKIzQtKZH0QiplDHcPg4
FDrnYyymMBl26ppBrEZEydomjlnzj8yKxwHovUH7mWgYpohppwqCByunAAR7TMzCqB7Z0ciAmkmG
30ZouKpV3+pw2et9XLZ4RF9QAVYkCNkVyeyLQ59fP6rOjOWMzrS0gpQWvLftpOveAqu5vI8r2N43
iwQBvvcVJrspnJ18tfkO0CwoDf0e3tcao3ILwKwmaOLjRXwokbLkrRYgQnpl6DnxcibtB4X7/80z
YMPv6F0/71JIf5KLx9e7oL0XemLaeqmKz+AuZmCU5Q1JAYFQWjef/Dtsh7YLJKCIf4/VAxtyU6rv
ZcSRHBXXuMu4BRIwmapU+i0XNZujbnnW+7/PimPrSLIFL5vGp1tBrCjz4Rn9VdcU3wAljI7pV6ju
oB+Usl96ioEhsGdYEquwMsTwGwkn08eCzh/dJexJP0bjTMb9ikYFaF25t1lEGMHsuXmoUVHdlwHU
qrweckWXOsctF+AfFeEc9OasB2D4CwcJqdiH6RohqVSiAajH66IRyQxYIU7VTI1VZWSNB0qydMFH
cuZ9J0+UtJZni0R93zTlwGOG2iNDUD7MYUXYLuciRjBwAyom19Fvjgky1i5qOfeUBUcaCh07EIEh
sgc5jQJ+uSX7IRxkAiHg0qitaI9hwagrEnUaD8BTPu4Npax8Lig2B5yyCiyhiExDAo1rncEAoPOv
lHZN+bfjnrTa6cRQaFUBhAJzXEFnZYHG+sBmj5gIeXHDsKLvsG8vA8lAxhvChlcL5pTRI60fBpGr
amD8d8k+JYnBaLNZHNlS2p3cvbueUo55FbpClsfO/emT7ifAJMhy+nJrKS4AwREz3NDmo8EIYHG0
lQ6z5JPD1hJAUJoxcoo5M+9poN/DacpmJ9bDjSKtzILu+JL2jAWZQn+zYArhM1ArPvHzehvxQW9G
P9G/ud27LGJfHiLLqPEI4kFR5YYufiyxfY0z/RvDjmTT2QofvXtxmVRmmTx4Iu6Pe99GjZWx9BHU
Hkm+iGrVSKzrHvJs8+mtf3DOTaqiQiGG92fOkgnfTt3vgv7eDphwAdhyvakHyp7kwc/EgFGHarxp
wQV13OffAYbBnMKJxwJONtCfu4Z940Ly0+w9lyix23DG0zmDWApYBOiK8ULlYozcnKT+gg1Scs93
LUQCQRBTZmhcE8usgNhlRfbNoktniHrsrpv+z9oXVLAkJi/9ipxWoCV76Z1oy4jn9KQgk/sMp9/E
1wCNF7kLsWjyNEHZEEzmyLpKjnjGoiBGAfQwKILhPIZeRaP7t05Tts7xbDHASkziiANhg/n3aLW/
lc6ObWJ5swe/qztg7IxMBaQ3+SZ0h21hx7+EkabwTCCcmoIktTZZzRe5Fiwy53nBhx9usR0MwsJt
VrjrxR7eE6yxkN7sOGeGJvam5bF+dcmciU6GdXQxHznWHXE3NUSMG6DM5qHNDgGBBUh5I5GAnJqM
C2+rpvxF3j6Txr335CeRyFJMa7PLhbT4LMp7+FEv0kopo8XferldbqUW1TbwFFeJtFjwHJ6Rd49w
yKbyX4IqV+qzE0spBVGN4gG1MDX551Ch7SkwcjwR52pgi4KUN2xwZfWO3bNJAZDjXhv8WdTlRLg8
a42j0V5FFZ57gZrOr09MeszKReqILHtsj7hKHqQhYf7o0WENyyRydEPa9lLaMhNJr8hwI60AojRO
js8EaNksjfgHZFFyzy2TVhwMR7JtxFJHINhqtVEuAzWOWeE7yX7KsLtv//I5ZBObZokeb0/XQABu
80oBnKF95zMjrjCNaK5Hb+U1T8UdlKSDXO23sIsYTQmR0buxbSb7Np3wN3OTIviDTcX1LSWAzOIr
fV634+f3rdBAdiWC9sRXhMdaZBM8xvDuPU53NMcEIVgbaRpBByJpbkF2qKMjpMhPOxIRLWkj2ky8
Gc2pq6ieGLT0IzLYb1ILQIHu+NcAnojOdvW++EbUYvM3Wqsy2jmQJRXYZYlUCtSSL/LApzkWDrQc
/HNcYlw/Cpa0xRdw/kVJM0kmrKDVeRfu8jdsA7wTuIUHnGYcvO5PmPUF23jvx0LCCtTiUZasMIV4
FdPeXSsoGJUBzgZC/sqxk76iG1q2p8tH5xc8wEQnckZUgifi7OKWVikAl8bATo9sBgFj1Z/COuQY
/hJ1veH9fCh065ODeDQuR+bGB+PnF76EltTSCxEEU6YZy14rYsa19SozteLYgPr3qLrGbu/eNL23
K/upe5TpvMxlUzXtAVq1N0AAMT3tnktj6wE0eS/Wye/hWkDHuhUpcXu6qN6yGxtePvpS9Xktl7GT
ekitv00P5f4LsJ2Ty2cJzu/iwQtCDFkoJhF6jJg4BaovLsb1yiCfrxiUxLVcrzD+yS44hfNKz/YQ
vx3xeEws5D87d8r54Zo7IE/wqJ5eSvg43B8E/KRtXJLD+4RXZyLR/mn8H4l6T5ajDWgVK/b9E6jB
KZxo4HhCPqvPuB7Fn3edJReiKwWZ0NO6uiQdALPBEwZMvlYjqX120z2T6wGFpPpdwOg0tHOz2pvV
mi7kldd6CU+khSJHl9h1hgcXcVuHDDf/hx4b+Mb9bb0GfirzKipSi6VunUOJt9BEPZVsu4npEsYh
ZCeQT0igMsNc1Xu2em7xpMhON0LyVZw7/DUsDidbLaB+IE/Oe0vfhlb1cTzOhlkGp9qs7yTeM/Bc
28SBhHBza0CM21qqH1u7sGWjkI2A0dYSjfR6w6tpYodYud1ildGAquPzSfp2n5ogLUobL5NMTlS6
p8/C5XN6RwCJaIkPRb7+Wx4rVRX624AizY+DMzjOAlPvtOY62ruEtt9liYwF6s8TDmatBiUXa3y/
/s92nNp1E4G1TnJnKVL7o1ordYVPmqLXB/h80FWPNC1TrC/zjEsX7uDIoICYoFQXqtOC2Artdjot
yHHU1g8YLvtap0AeYDfier9yipNXZwXDqsn1hx9rmrLC6ZMUXeCWz1zGdPhzHV1dOPFh4g7jtgx+
7tQ08iOen8DYVbV8P1a7HXRp34czFksh36Af3+vPmL2jDtUHRD3ZviIu9KiHQ4kKwVXSz9AO6+zb
9bilxVx5oWzrdrJbVN30sa7wEUOIxAPcHmOCPucuIBHxUd4XczEgf1M+pY6BvwQYsZi9hn1ZcGoo
ooZ0PBYYgRaf0t2hcD+DHA3bmGoYXOjqyfKnJzf63cd9cnHo2Z3ittOwO8SScJNEa9BBJM/kw9xA
EjupaYyHLxVN+51Yjq7JTSACuUYYw2ipKGfbsGhpWPuVW+6WfhoU9ZzOnqHXV4RlMl509FD8wnm9
W/yNMbB0ZeUOjInVodT/HsD2nCgheXFM3MMtYLZl2WE8MVL/r53XswcfC4OnHQNCadCWV6ICmoJr
ppsPQs0438Ho+vmGqGM/fOFe5np4IwERUdPfyHZnHyfb/EoxthH7cu82cnnUaRhn1/G+2SV977lN
XF9MHs60QsVWBuh3xU2SlgIJAkschfKmO5gRkXR7LtRRkY/2FRIKv9wuVLPHpoKf5qFUM+ctqIgt
uWJ7TrkP2fsKsVHYJ/7fjGuY9g+RP5GLc038038i4fw3ip8p67iqjYC8qQxaQYHGPwF30NtXHAYN
wbtmLCE1wkvC9Yqqt3rAu46F36/+50kJD6T440o5hl0xieVitfZodYTDrDuwdpyiCGHyCtiJpfD/
cT2wBQSwaEwor9aEp9XUxSmNXi4snzwSvT0t8AdUhAOh+0nEo7MJGTl8pf8wM98y67LhAnKbf6RD
yXI81S3pMZEuyYNPO8kEkI3SdHujQVZhT3b3I5dVRcKkDrKIh5d3ReluvGXkG8IUdCKP4YlMuHfY
dquNb/3DSepMXZ2Iwwe2SDtFecipCHquZtTu+6w4fDQ7mM325/SJX2Oi82A1NSG1fkeJdoQ7aZlZ
qBbJ96pijFdCLTxf9z+zdF00GF4j9j1rjCO0cViuhm3+QVxrqKuv5KxelTSvBhI7YObgIuDhMUwf
HNX9092JwVAN71lsXpITdVx0+pCeq30ti1PfJM+RywHstWGbjLhdNWSokJiuFrcobhm3h++kA/Wu
71oySvmyC3GXe5bR/1rpBu3sGEBptaQknkFePt5karoYq+uhE/ootzAvdY3FwP05XWoqiW0Un+Q/
fs87yPb1bJ2O90tHA7KGOdZ3JiOYCS2IsR4/cP7brT8+Rnsfk965v7PXOQZXDnyx8xMKXJQiJ23F
do1ECgs8OTZRTLow4WeO4papX1G/wp8AaozhAH67FDTDprSqRL//Sv2F5uWddFdLX+tEkenuUGok
ZX+sIPeNSgJunI3vjSfqki8CtAI1QuElXv0MX+0WxKMWwWAIJThtb0sHjewrf3EluZcWYMfUvDMF
wHPXI1zvgkz3xagQgon3fXpw6Xk4yRJ1ijK+jNINJBVFxsv/u7rEY2eovkbUa0Eeree7AvCNvmUb
2pOkqeyoQ/dEjqKlxXqvaTx8A67f4KVxNrEU3kAvaDtIfAlw/p0kJsq7VnT3q03HMGaBGRHXIGGt
Mqz5tYSOPwfxdEnwOq0fdMiIdun4Wz5m8HxYEE4EinN3rXqMPqQflj9haXhaO5mQB/fqHhyqGjqr
zRBYEIg6tpFVOxpajGh0U2XI6JbTl+1gwoD+TvE5jc191GdGiOJ5zMwYHvKj1cyagQo7QBcHvKP9
1qM1jewBp9XHO0KPs4rHF7XG6lH7J71eMe+ulc4w9JCJMJXJ5xK/LMsDCGFM7a5nNXehRyiAkXPq
tHtme6MsfGtFAgQfVIdoVM39fd/DMwgkoM+71DHQiI3TjPtGZg1HY6RC1UjeeX5ARlTjIcQi+UYy
Z4Y32NmRYOeNB0qJND24y0hNA/iHeAt2QjLFZXHFxxDKlyImLj7klOJQ3wBitQLPWSxsshYrO5aK
o9BhhfaJibPTsTg2U+jy7m+VP+vye2zb2O0b5wUGNsXXiazhxKkVaW55dyctJFiueZTBMZ9qBvOR
34Y80sfekMjo78hvRTwyLpsfFJM8HZNNCwMufMLSuD1CcAMDnyMRGDgLdjUCA3bYnAn5e2axJ3j4
Gh1AxQ9X0cxAH5588NrB9a4rYK3SpwiICMJefdJK6xahnbjyhV46jxyODCFG1PPb7eakA8gcud6r
DiiGP7hGVgEDyj+kWvU1WaXGV6JcwQSUd4CyoY5/ME9Hvn5RTACaE84FLH3y+72C1izdLA7g/xlf
LSmkAvB1aLfpAYl9/z0B1k37C9gN2hXT6ZXJDLLpVkyx3XMQ+5OdDh0EeJqopRCZk+45R+2wKCDy
eMgQfrguGedT1WeGxLiMveRU4FKsZ97CVNt5b24KtvOKbcW4vV8BIHPEMSLpOn3R2d45m8ocrqdV
DADRXlxWHr96cL0jD50UuDTXYjLylCbleyQLSKJ3htYWmarLQ9yDOF1WEt0lrsPR5gYVwzsY9DmY
NFmdMZJH5ioc4YsDpBw2aEMrw0/fMQ8tvuZSo3iSbJUYxRt3xUc7QKGBjn73SkjrBh22WErwEv9w
lyKnpucOQx44daKyOlO3UbwOGhUi2r1W3uwZyBxitmSyUTOu562GOW+jSb0meLNtLr91WpmDyemz
Dz16qnHwmTekaX8/awTK4IpcKidjcqjWmFwpWGejLQeACkEQhfnIdp1vzQWHZxJJ7xfDuYxAk1kO
xm53L0heQweoF1TB69k7Y6kKjxoDH2lkn9iPUbnXWr2yBmcSZVL1uWtRIogHXcU/EDUkX2gJLl0v
v99SiU1IO0d1CSbSV2+qLBN3vqGSQOKH9nIAzz0FazAASuqaTmeh6HUAggpVkUGxcBMy9H9KDKu1
Dk3IUL+G+OJvKS8Jxl5vhlRMOy46bxy9KhwemloEvRQ04QTVwVV1FTWchyNUwKS7yPo9piWhOBig
P70L2FjDpJPGGFXZsjHbOi3IRE30A4wYHl3yhzUREzBfHlX4NOl3C3pmE4t4Yz0tmtloC1mXXek0
G0zwNm7j5aE7wQjceSzBJUgR6qJQy0+XBbku99Q21WQiO1K5IPwu64mMlcPaWnAl/5cfiTN1KrNm
Y4rA3dp0hnTDtk2dbZTa4qLaHFKy39C8YiZlo0z3UR3SzEU7DOJUNpuKVigMX4Ffd8X3Lipv5HZK
5Va7ja3V1GNizd0M/VCGzCTFBPAfKVWtYZCcuKS16c85J5ivPaHwImwV2eTMNACrEcJ115L0Azjl
ahLdp+YXC42LeKU0aRKBtJydZYq3Axneu4bbDGZyrt6tw2/IvlBFt5n0Rba7k6ADUKa1D4YTPK4/
H1OH/LNEm6q+7VmN7w2ERDMQE4hhIpMypXhRbq26EF3Bg8m85KBb1PE55kad2+GwFptKbcEZuxGG
TAcVDcrkHstAtrL18X/T9H0Uq0jgq3cinT+byvlKOC2RktD5z7dP6gA84o2LwHCc8DRNTd1FjkCf
vA2nY6vVQflWDuYzIl6GlFnapwoZKa+ndN+Svd6bFj7FSubu12/8IjY7z9p/0yqgNYY/0xQwfEyt
6QeggIydExHP7CFGCMlvneDXrhIeJw3d1Yj0pzO0BGG9Hp+Ke7x09fi4dKR+dJtxcCj89NvwHAW0
8fNmjj67m2MHCG5WKnyIbVkSduly7kQHtZMO1EPkTtVr5RLXdGnKhDrjELrpjjIXxaS6U44GRu7/
nhg7KFX08tFcumPW7UeIKFmQckllk+S7UZ4W0tKvfDkAu2fPV5N73qiNOHdhxP0T7sYk9hNVCsyq
7nzJyiTQou0zMwvVi8omPBt+nvVxPVEYqS2KYu8FX1ZvpgQ5C7vDAFVlK9mtLoB9FFe3HjmejnhD
09pRssCsXBqWa3L45B8RB7v5G7XSiIeon8Wtb7BuCX4kyDzshabNkEsCNawIFTFO/9r2LONjqHJm
mDzhxyicCSPObuJUfCTQg3x2XD/b4FHf3vXKe+gXwTfCWUmmZ6iJrJPpd/Sb8l49Oynw5WKWlH7V
EjOije0689Mm9Qp9Y43J+OxZaKBT8xjR96Uxx7RBwVQlgJaw4+irON3DBWEBk+Q5q4eH8+7wSlvH
z3SX+j0D/aJrVF5pY854Ajew9Hs9JfRzPH+XQgDsGkJrzEVRW88dF4SsX0KDqUopBh6JOMV9GBGj
rRsjJcqOTarv+PVguKlV2SDsEz2OfJ5MCO43gUwHY9kvp2WQPK2d4HWjgwnPiQEPLGS0NQb3uNUB
z2gOOQukHmjaLHAurIBqpAbU7ksAD4a1NlYkjT+1UeTnxsbwq/eUwp7hox8hPhhDHEHTlnsPgIb9
VW1fu6OrsVn4oovB15E5rtgw6mVUSmuMheMJBjKd08Br8e7/uRWnA4x6wRNflJ7rMC6K132wPqKA
6f93KE4WK51wc9XT0F8Qj1IIXRIH5ILj1OXKcM0FuteWb/g4omC0H4soGiPZ6rUZOp2Iu/3Z54Ju
ENdah74AGwNkxDaONtRgZEmR5LdaDWN9LpoydjcG7/Z/yAyhWjlA/pGZXI3BawxsxO47sCHjg/gc
KaOdyf1+X/MgIcEd8JFufnX577bcBVbNq1OI7uU/2WwAFTaSPmHjXPpuyNY+qySMO3iCDUxbj6j9
buVhKJMiFnVM9WOXkkiPyvCwZv2gFYMgbQH72dcz6/F+McXQx52Wex23QUWsE8r11gDeyGn+gqZX
gp9wJxt1mztgW5IHFNQ2tKWEdwIkSn+2o3bw/uQcz9ZTRlFJy7az0zknn9/ZBvZ6uTGI6EycyYMg
FZL60uNrAw6Ja4j9AN/LQzy+YRIPpAztCZe4N68L4H+VIOF6w6PYzNXmqWclqQr5W70O9KS7ZGBr
+uDm3EtXCUt90OTcknpexAkQBI1xjasm0p23eoQmmlWbZ4fKnCcwpVr2EXlq57FBig3xEhgdqgz8
VIOAkvKWixoibjIIY1gIlvv1EY+iUOj000hvmY9w//UE3wOQPxkDt0tGAV1+M6kThDN5sS+cyxe6
NneBGR5N+wMGNz6QtsehiaLyHb7JLeZaFAiXlCQtm4cNO0v/jw2lXWJ6srVarX3+lS/sH0MRkX4X
kYawulNyfSiVcgXeLI/gTDhL5oJUs0FXgudFPuVzkmQRUEFi1VZf7ffOkxmn4dP//U+0ba8XbVgo
cyRr6R+kC3/MciaIqCW2olgcsbAPyklS8tkz6SsBdyYSMAMlCkZY/nWInitFah0iFRxYPbwT6F5C
15iu+suYnRxv7Jh78mQtVhNFsYw4d1CvwvRP7yZ0/NSkO4Gr9tfmDyB14PO/Awpc+oWMKJNGD6be
14qS6q8BVdKQ1Q21bPTIqOX2jm6l37EalS1vVnmXCohOgPZpzT6hxzbFsUqu3E10+rjs+C0/evnn
8FMf+J2kIgekVk9NNqlWsE578jrjs4RvlzWDt3hZz6TMyqQlFVAglLQHebuh15YUdZwLcp2u2t/W
j/63xpuR2gFS6HnhXjw7ybpckUsg18O8jsIJeXLHhz5R4Sm1Wodbht4rXRV+TtPPDHFgNyK4GjFd
ws8voO/uYs44/t4lDZbX71s8aluPrdBE8ZaUB0XWRhkN0Zw/ULvPlBfVBEGIt/2TYy3l2v0AH3OH
s3kNkhLmykv3DaeiTVWaiW948Ws0ZH7UUx/u5rGty2n34yNA+xBllDnhznp6+yu5CG6hmFjsKvB2
dLLP6fS5qlhaHas/7/mg5A7Af61YfzjT04qwg3BiOkfyfYVfIF8EXn4s9zUP7yyaP2KbyDddQAZb
iwlIDLD46Z+9EYBcwY0NsiNXR77ecM40Rw8r2FgZdy29UwS09J4xTKer7KDDbqVI4o2yI+iIHl7G
Vve15xrS2aPAEgb+uxDF+7itXdBrKsxaZgbQ+7B/RwL+fvj/g+7veIbKJEfmLiUAVzh4n3QA43ht
DRg/MmKUWi7Z9NZPRlZ5jIdKBnqyrFL0yjEcxR+t7YplzZ++GXRslI4/j70YWuPYw03aFq60sfuF
x3M3VcTf7SoxxfGrNkvQSgTJ6WMrrMlURU7DWezY/M4g5MXTpIyU80V5n1du9e1DojWw4/IfqMws
dkbKx6zM5iyDfF4ng6oa9PpL/EM0xxSyL5lTmwjVzxmx5kjpLCL6TZ20JVeRgY1noVbmeZPhrR3v
zfcM8EfTVeRpMDkIZje4qlDwvn8ixxPqcROy2+n3Hgxep5nXmF0ZIhl6sgqC9fXewXYWULAlSTFo
EcorwuFT2AAOMx7m06G9NEw165iK/RPt1Nr78YGGmv7KwaJksYXQkOIGZxPeYjfG8NiS0ihN8Oiy
s/TPDLg1hnvNiQf78BU9dfn51jhH1z+Zh9nNTEflCWSOuswGNrH24PF+G1zi0qqCeJmf38mRf7EI
NjvWTY1hUjS4JpkDvw918UM0TCbZ6mzoLvUsVDRaDnZ/xDYv+i0KOBWMSjjZsYXseCpf4GA+LeUv
IU8olTO+I+x2caDHhRBWvtN9IusBvYDTUcAjEuQt2SG4Kes+dcZWdoDZ/uZTB0D3rqjl1rc5tHD9
Umj7wULjNn/hUZ1wRx1yuX5EBT463aVFSZbvEDJuEuie75IE5zLXR0Z5aWgo+u4ndRLY6JORttdl
rSaKmsI8p8MnEYcE4ipk4fqQq5L18nINqc+w8Fik6hG7fqnK2wtyIxwgtOxbbwXzCD5OaImA+50V
qRfgZ5rzWVcizBK9q7FNssr3uO3H6p69X4xiWfMTNzirlZNVhrSlygpe5KmcJjOLH/xRZyD+KDBJ
VSABJjkFfUvHufr8ohlb1P28Uy+a37vrfNvPoiW6GcRllNtu/9Jx9Mbq0rJzZH5B8mhpMqYkvasP
Q7TlTG9OoM6T5uKdg6eulaXtZzAlvRCUdVgKk9tzd46gfuhQAOZWs6Hz1Ga+WdYY1Egh36x5C+vr
34b/ETyGfOsR4sZBoup4zWZE/lD7C3RjugDj9ZTCXVU/Fymj0B9Tw1dl+IWuNHoWyIFIfKMAlXzG
Q4P7AI9MW7QOj0RqKLlJAOu2O0+c7oyBabJ+nS56nUw6Mz2SnvzFI1nq6JY4vL4yoMh3KlEBqCw6
9gKlR4qVlF/IIDf/QHUeVkZ9gsHLg8BYLW++LERbK3Hr1wW22OHEb5g6kZ3dwB0Ym+I2hfHjJLCj
y8X2Ys4FQ1vgl1pss/mKokf6SrNAfjk6b1BsauNXAZJzmZewmvgr/Fsr8Dpz+Tb9KdXe5RWCupy/
oteJJHgqZ2q0ZbD2GLU4lk2D70LnVaF1qrAKk6+75po/7EJZwkdEnz5xcfvjJ4S+UK2lxcs7u9Dv
SJI4qMnD3l5lDeu5fKD0a+gUN3cURmgAqGZemjrFxUOrW4Yq0yqCAqf9MUn07r6qZMxhOjl/m8pb
t+lLtTlH/B3WJ9UqcNnAq++J3tASJLGXbjPze4gzXXljZKjQSZbZt0kklrLh2SyzjXmF/EbX1mgL
SGM28KSLYWyil72p0+wHljyrnlzRcdU0b5pn6PeFhJLZbbz60HPwEKcSt9MpNMTnL1TjLBa8WXk9
sdqMwIAlxukOZapcgGqSOoB9pIA9CsWFYzMxqFdOXG+W8Rm+ieC1mT31AvNZRumk9WayvPauk2Ca
MP9cFVp71mdEbZNA2Odrim2kz0Wue6VCENWg8tCzmnAnY9hsPE7lxEwsXZoWISxJeAGK/0O/mD9w
8Rq26T9Njp7c0CxNKvwvo6USZSc3uxx9EOBmTj8nypzVzWZzeEvFvPy1/KOrtDzhTb/v9j5Mliiq
ALwlVTYVBzkCd4mcChimGxxqGKZ0YndCZb5znIHC2CaZLY032cV+f7hl+fU/Dsls4/ma8AXyJSeT
DVfjIm+AaySYf0Y3HBaqsMbTXeC1saNLr4xOzYewIad9gdW6KyH6ZpO0xfbwSUMmWchqO347ymOl
HJwkIfHMs2a/JGjPptmtewCcmHrwioVYcMjDCCBwl1zB6aj4pXfV0qjK86olMtOxFffNst4s81cC
V2831xVLmGiJX8iMwRBqpY+AQzVdv3uIBIt220rx9+ysYwFgiSGls5hVHso1oB+H7xK7TEyWHdqV
4wRbAmUF34Si1c5xjkUnAdlZzPU3fxznI0+WbMZX/tJxL9ZgyK4AY9nzJ5L4TEzCnyeBYgdBOQd/
cBZHefkexgsxL/xwqM/FvOlB2Ct7bHDLywhfpyc+m+E4ERXn1bViZ3l6eP7j1iJ5Wu9ttE8ZRTYQ
vhPWGSlMW/9Pivno8+LIPR7izqE1hUGhGT6my7RN03m3Y1pSEkGwGrEYICBmgutUplT6BmhHOuXC
kU5QgFpGeqGZMbooVgYPqolmRgTVfjKbGIzVIwLxe2F7QdA8xDkBTa4PWwPldu6Rpk/Fg7FkRRFy
cVpSzwiUiuLhuUgtWSfnNHnst9NPSDGrWfAxbmLGNm2MJQWtk6gO7kIiBPemBpHe+y9LrwaoB8J9
w2srXm186mBjuoKyM2zKFVtCP/ncA4HXP66OUBLSr4XoV2xKJVBa+yMvFknDQa7K9/w2wYsXKcoY
Sm2ATYtWjcqfjxe2OH56hy33gWWL3rDdBdvuOn7r6JEvS7CGBoPyBXGhWT4ZNpWvkm0oGvtkvo3b
+0Y0uJlNi8DLNWuD1SJ80/Guk1OF+kqJvpeure00acaf+E9uspE8qKnMnpaLEv1RdZCMY0g2uimV
mG5drEGvblOfKnZzo3wXI5AvUFDbxF4zjDcfrymuNttmPQNiIvtyk6Rkdx3kBPCbR1Sq16Nwrrgj
zfx1Mpn8qqdcsQVgo+t7AFrwEIQKtvDJpWOSbdbZus5H2hakGPpbSoe+fmsNXfjmBT7sBWtkrshP
ieZQJKJMukCynQVl02iXYuaKBpYIdP4v29rt6rPwv610ZOxq3fj+34RPzJsbNynCoaHYNXeB+pkF
D0U1yQ8EswavSNzn6YViCxjkiy+xUuQzTWuKjl/cSAjkxx8qllnDMBtBSNOFNpYbmdPlngSv4h2L
EP582B4OTA9L73+y2JJDl6pAEeepSEqTZKyXKpsVVQhRFEKsaKZbjuUeR0Cyk3sYADoY9Th8L28c
A9JC3CFUuq1BBW51vDJuom1jJbOECBaN8QO3sBax13e/mwOejom4fBfR2gvAntZFp4wW7uSuMYbu
V2IdVH/6ch0MAddGdbPivxvMgvN5eNHH8DH78KYxwcTkbzedyc2Mv16BXZD2vMkZuSpllvyL5y46
nvPinroUshhtfUBZ5/9ZAOVuB7oEmiVFu5w4JYSv37Gi617S0AiQuIZ6RznHRaOGXLSNB0UCfEdy
pvmH3S0ME37H9fn11B0ExUKIoWkV8ez2Vsmn1lcxnOPc1BZyizUVjE3QEuRfsKf3eYZQGuQVk+fA
cJ4qli1ufTFsGehXLUo5jyBg4FcYNC2ZdwLR/+59Y53oF9PDtzGuwinVko/QGgPt8eKFuOh9W2XA
Qkge1PwQpdKUH+stGV+pC7wv7r6dfrNkQEUJyGh1Vt/aWBeMYbnnquFmSP8RblN0EEBswP8pZ4qG
6CocPMkUv2ouD/r924mSjVETeNWKhsIOVMfBvuFlHncEElNincIEjwO/94AmeqrznCyF9g0KD28R
4JxhsU124zjrOPmpye7zq1eHZMam56/rKugxLPKChXbfS2jaE0LFKvE5a99xycZQttudhNpCeWye
YKEFWf5WRKAPMAl5ohT6b6Em8JUCwwDtCZZrN+qhVpPN+rvQ2rGBVOUaFK6TKzMEQhGFLUNZ/iIJ
tcMOgDSIu87pzIfT48Ba4rue/DFBJ10QwiXJVDLJzJDon1mxDtm9Hn9Kuumpg59QDR2BUx+PeJ18
Ewo8jhURXmmK/BUh2MxIMrm3Sndl76LLxPC/gs0lmBgOLNz8fSTYieyPTdd3ov8134NYcJJnEO6Z
iV0jRy2GLxKhoRJQQxaxOjfYmq5qedg4hWxj9iK1RD8Y0QSEox73HDqJ+LtTtbXef+Pv8gD8iW0U
CT7GDFSfrRcAoWJ2Ko1/tbsIh0U4pA3W4nq2dpW+9aPd1RPrWzpKbFxt3oM/tgtFEV4In9GrKcwM
gV13P8laar0LAmogRowWaDm8Zt6Uo7N9lpOaS5OFZ6l78JpF6B7sSvjr0FeQrURUaEGGzaplV9fk
GxfULvPC3J+ewyEd0ivOpaY8k4tjk8UaNfypsmiB+cCg3Yh6aZYXlwYnoPLOCsHPmK1eC79SZ+ix
v9iDQhtOf+r4E7a0iKglXbgM6NwDUBcuqdHb5EFmaF05YTul4MdijEqYOub9K0poUeZiFeVrama/
TD7OKENL7sF+cqgxeYULjkxLbrVmucBvrvkfJonFhno4upc1CJo8L1NRx8tzyWv//4nZch671eCh
Ow8Z27lNPLz0QlTZt3hHw08OUL3rtzBE/+sN0BHQhNDq1+Bs9iqzi4kzLeMszPEVlkiORIqZJWM9
HziEcnK2wANgxggVZYjzu2xlSkd7Fh33ZUfiYrWP1zPkHF3x63Ktt+MAzVG/1rLgBcimQA2VHFSG
IjdNlRZzeg+UCPc/Eu4PQAvO005n2w8V2PVbCPlv1oYswkMRvT5IUqd7fYtyL3eoXS8uv3VWcUtN
8HoZdDRNwqBsR45wvJeYfuEZ5ebfRr7ljgL7qxFtesKSBZDID4C7/B0/EshX19pDI8dnxPa6qjBh
tC7oC8L1DNBuHAb/FvZIJqG65RXoCbE+XPt5UOWbNGDm+gZw9Wuap+oiEBd35KlUoHNE89Vm9U1X
UptwVyNZtM8LwvtIp2YJuXwPyqweo/7sbMFlkv7KPArfYgdfZGCjPJk3srG3ncSlLPEk1/jghRs+
EYQG+JY4kFDqsSKQbQtfM+HQZJEg2llMnz1ZxfRaGrn65vYpljBMJLfPtxpjGndLUekVQtvaFb6o
bZjJbqWvxIB+wfFxfyMwEIIpAwmLoTU2l575n7/WD5YO8S6O01YXUSz3tY+8hPsIzd+ZwfGOtTgM
ZAB5hT1++/cjbe72NwzINB92y7mPCPv9hxGzYLPn9dFZiWJ9sX0oJvDBmEb3AVKmbkEXCKIftoh5
8bqSbiJLbu85DsOT8PNi3THLdA1bDGn1G6NGbVh+UmDRimIPsAhzMX9u1Tur3Vtn8uDNYqg/cMGg
e+RdFYPLuE+Gdb7s6nnD/p53xqkf6z+jWzfjz02hMabifttdewKMN8C7LePlr1R6zkQVxfObmKCb
Tj2+tSKWjLu1MqKFdn7lvySPkei9lO5iYD9hD7Svqe/aZyYnakzx+ySEvCIxGcQ/bl+oV46aQyIw
pkr+Qu5L1o8PhEaIPmSEUGg6ZTt1uwqvw49hppfEtwQ00jGB/cbr1o50z0hAMP7r6nfKqrxFahPA
8Vgal+B5bnJoBCbY6xYGqIAwM43zI7IYz/3b4+dGGjEu0ltECSl17jVX4KzbadXN43JlDNttUcEY
KZ7ncuVnbc1FTGRdXjWP7Pd0R31Ma6A6iVttm1h6ICcfIlwDnIHXT/FZCXM1qepZPgp4Pb59icI/
Zp0iNkTIdy3+YIXbg7O6QJt/jx+5MUDE/5PgWA9MhKYp4FZhn8VRqgxuELGemoUPY1UH/5wAchlW
ve5sOMgvzIf/cwRrwv3yJKBTK7sMnCvXMAaFCBgqsrlBRU+6P16uo5l6aVE0geS8eKJrd74Z0A3g
TgFwqb40qrsM4QZRfB8lzXz9QnBLDEny7FpVMIbR42MfOJRIHu+OMHz+gyYr4ZS8yV4cImwhc2Bw
VnDKmisGr+MlmPFhZcMKi79jdpPFSkyh8rRvzYUIpULeq96c3sUXEFevPyi9Y5I/NypYliv7tcr2
v0vUIBtpt3EmK9E3hffJbRlYblXZtHC6KHeb5ihhhYAcmUGn91if23tA1HkLqST3BFujiJWYuVBY
+qXH21bIfY62lSyh2NHoaU+XRNFLHcN6pR/hQXZOOJ2OJKHxazrgWg4KfM+E95p/VCuj/nmi+jdc
8P/z3+iTLJGRfnE5IyJUAIva6ixp5AsHOhZeHInQglQb8UT7ah/34iScysMjSUo7sYGI4Zro01yy
s4PnFRaXpB1T1ksBbh7+cwRSoBMdKdY0nvYWcv6mIyiKYL6JU4VlqmkcEKmpFcUthXdZQIJ15/9+
arIPX40s4TDnZ8bw0fZTF7LdADqSaJL/zL+rvX37ZTrzcwshrAENtl56ff+WjNygQA+G3pFAt9hy
fqiLeIHNYmH+//Q198m61rvL0l9yUaFmAH6+Xxx7gN2kWlTcP7ge+K4311LEFTyQmEMCLJFNFr2r
u6KFG27NbCsR8y/dUM+FnFf6ozIql5ZmvalvtqNC1/tEWT6+aHKuRg7ym1XC1qWyFUOOVEbOqYeg
oa76lGQTnaTaIIADjzi7//w86YvAThVmqSvGMB22I0u9SW9OJCS5ugD5FKM9J5uSzgcs95bRqfGx
xU7d/qyvdUnuTzRdwUXPk3y89MzsPiigm2N5lFM8racwdyPmtn3l1Jv+urMa1AsxEgS3J8Si+unT
UxtkQzNrpWLJRqbmKty7m6WTzP6KZR66BMqiTyRgZgvz/g7orI37T265nPReaYJg8CtjqvhE9e3y
pEu2NZbjytWIU3vxm6Ny5iyAaBc9VdEKdSfLVtj0KdB2VHmgN3HMdnYZwDvcRv1W7aXyrZZBL4NF
PPewD4gvBv1v8O5Y0a9OmOpyUnev5+fvViXMX8sVh3xVHJZCIDLvaPP42wKi4RFMG/vVBEMrzcTL
WfbqHthFPP7EoVOeJ8A7AriSFWs3hbxuRG1ZOAxHw2RhAAbScVUv9Lrl82n49gCL+lMmGgQhLMlA
EaZnEvp/0ZBaxb85cIEKTh4BLuuGNanDWgGsLOq9+zO7HcuvVbINnEcdps3pkzkkKsKuywNLKsEN
lYWjjs0X61Z3nmqWjSkZ6hoaMj3jF5spt8bth5Eqc4aF4vGHZTp4yxA066kLT+3ngnb3kbxMeOMD
L1TuLcQxxrSEF/L8CPRgMlxjm4LAMLaBBwyua5/CT7yqunhyDIcD8r0eIOinzjo5eMtdIaC5XySx
aYNbNCVP0zbTRx7ZbzcIJkwFuRovUzIaF85XhZIhtV/4BlJiEZmp8F6CAkiKMIXGyaifjTIg5yXr
tttlyQMg2BEJLJLra8RA8bu50SyE66uQEeJHc9lkRNuBi6jLDnkL8kyJZF4wHX3ysYnu+Eh1T3yu
kXyLkC7ni0wTJ+DToHgQ2p/KDV58AToeLhYurGdZU2nklJKSN+uSBsIj3Mkscba7E8l6k8XPZ0RJ
6EPpOi/pnjkfqBLBnIiQYbgKi53bmceERVN25rYpO7YjRVl1e8vJv3rPhQGXrXT2OPLfkyzTAFu6
fEr57g6a04mNlNW9PdtJgQiKbffUq24fS9lk33TDJs7vsuroo64TPrWlQhC92q2mGX3UJ29zVtEr
sH+zLsu3ALRObqiCV/Qd5ett/iDrIgWW7DJEQfMVqjuvtRay06iVbkaAl+fCgarDXqZBCSLD+iIs
lArsGZBiFVHLJ+ZPNWQFSEisogcynACNJNM5rwCsFh1UfHurlLuN4i9dUBUMi09AcklTcfuqt2nF
yQFYfXqoXlEsYGdFYUgsIGGydT9AayZ373Uq6H2g8tgXQH10yP/6uWPlzkXGs9MjSjEVaM4Hk/G0
1voFH7CJcfpxDQ63OgsycmYeTPCgOZTBNMa2OWUaSROckz5b/sWxdY1rc2yddEgJhOWTn36wFgC6
t+ofb5W/hErvbQg4oaf5zFhApQI5P2QJEFBj67mX83J8KbCU5MuwwXMxtpzrHKs5t7ud9b30Eo+Z
/fvALk0mFmo2cGc/7oIQCWGs2xc8+5ikPu1boc6mUl+lkB1KASne3fSRHpdzxWbybZ1zQ3uDRowC
Fysa8oq+mR5jxNSjXaHqo2CJWVVyfkX6SADtTQ60u9c0lOJvSruR9KewW91DMfrNZoXwejVuPRja
RqHFwfChMFuDaFlCfIA0ZSkM2S8vWDlPEoUvKMHKn0Ql9perhObJvPD4wuF98VFk21ICGvKr/RKb
iNwNSJzR11WCSLncV3favLeqxvWLXnVrNc1sy8+ErtMGkZyyPb52x1rI8C/pfQzu+NaO9DpL36vP
CGnV60qxBsND36XmnYlQq8/DoEagnkrg5OTbQPYWpCuc1k7MshI45bicOOyVEVhQC2OT0gf/c4Fh
ufd1fjGQWtuleKa4TR4PMFsTj0XfttwGNTINyosZMdpb3i8dyGOWmoKk3d+DC3s76X2R4uMZBdb8
y1zk+P2R0PfZxr989Os1b61SC5SFNRbY5RX7C+Z0R0UowEezRwkFrgXHR/1aLgNJxpNnAopvD+N/
P18VKr9AMJupi1NXhG6SZeBKiYZO8u0GG8igXBfElyi68hXXcoXQwZUEgb8fC7Jb9U54W7/sFTTc
Nzm4n22IOaye0dQufU19tSEBB0eXCYx/MuO0EHBommX62FNw4EZrSnR/4msVzwvI2+gOTBAIQFjI
RiimPcaZ/hyDzIF3ez/gCLE1QSVQrgNxtqBzRnJqqNwhUJqXuwQOgJaQFG1Wvw+4Mory7XFqXTBq
nfLb7IkbRxfUjk8kMRaY8QGp7++FRLU/QC2acHxAb+yhLTT/GdVA/vWEkN5YBqPziQFOB+GYbFis
8L8Vn/9vkvTOmLULYW/DK+uJkG7oz/AxFIyJbvEnAacbl4XVFa5yrme+Wp47MkukZHnBh8G3DBMZ
zftatmQpAchk4hdLpbbNil3Lw7kxv/bXoA8vfhRQF+hRAU47HrDyPmnKRqjKzI7wd32n+0bnvlNI
AqRK5F1OzU9clWbIfR/Pn0WjduBTa8b/u7g9K2U5baIqqND2/g3snnsyR/2zOsDufZh5oz4VfdOJ
ZXk9Z80MddgbXmnyIsvPG0aAaxLZiwDRUvPFvR4Y37X1e8HZ3r0gEdP2kIpWQgDm36VNsLOqFYI+
Ugx1xxibKVjLALD3wIHs66yiBXnZlsR5lI0FVICEJx8YYWsCnZS67LKJ7IiNoej4Nh9rwzMEPR7Z
nGT5LzmSC0404kxYEnidsGfoZMwUuhjrUFZvF9YzCK6AcgmAR2LpaLC5ReuLJTwk325Di6C7nz+s
TRtGuawFxno7OPjy1FbEk7L12qtXEosWXJw/Gf+bqU4G4H5A0dK7Jl62PQt2l72sERWKKgiQEfou
dOWbNss5PemTruxFuDvqRS1QHZR+PemQKkmt5tZ+n2/ZTsL4sQB+yx5NjuHMmgg1Z1qSd21RHNT7
gCJYoldWLt+zcSjMYujMJFg5JCj8+rHLJfqHPhtaEMd1ZZv630WvpI0FlmtQzw0X8X3YQPqWAtrj
SRCnOS/dH8c6hzYrWV9j7/2vMi76gbw4V60dTmk1bzHPodpJ75t5tkUynn7nilodRD68jaKbPVU9
9lOn+gtUhXsTEEmH0Sqqd+qBU+/bxZuzPNr8leQO7qPOC4V38NUO6gR85x/bzoBQiitXWvrAEFmf
gC5ywLRn7wdMrJD2nrs9a2K4cHDFB9YstOX1Nir56tlHmpLgKH3LDMsjadUEufti5K/tubf5W2LT
pkZa0DNVguwEtGf75P70RMxiyrPOgdi8q4phgniqTY1mfo2Xg+Tsv1M215lVNFZbXL+0Vu7Il1P1
gyqnmw5MkzoQDJikbGixMwQGquGYRjby5J8V3TJmKrqUtYaYxJv7GROgCRRioCZq8ihUds8x6FoT
tjHeOhKPkJyEmaCpbCgAqaewQ79bJkIi9S3eP1zdhGqg31mKLmYcp6y2TXp7Aa+2EyEGtQekGkZ5
58YdXGgdFSmd9FpW7S/Qzkp78DFVb0VafC7/th4iY3efO4RwR9crjZCX+S5AL9CoQlEQuYn0XKVj
9WYdujxeLFpjjxMwzrxuhuInH72CTV0fg3dtEmlVio65C1qLt343umsD3AF94JtBlpZ7KyPZYjnj
2h88v4rzlQKW8K4C2lWvpPwsMHLNqqFHAQnWLheUj7Dq1cjeJPc3ka2iIqR2i5L//e+OETGFjeaU
EiWQ6W/wQJRX3ugV7dRecVMilvTAsyfVmUtILc/5j3VbOQysWZFJ7UFbc3COMlJVNfMyBRHrXWeJ
wuFigNIygDBBjZaNJQs6enhCc0P0b825QJGq4M0HEuHGT4tFfdupv69FVHOok78f3xkPPpG1hCJ6
H6+c3ikpHEAQrIvZMiTYKc3PLfkh++1PM8A/uWgjVaC4FmuuZ24VvvHjqrSexjlnSaGPbVKHgsJ9
0lyagcCTBzxNcNu4/bffGEYSTW/IRKQwHOY3kOYtg9E/CNYMF7gEhPyqxRjr+lGTMXUFYrvhMqil
24dZJtl92Lrn73f40qhLFIWRihoMCBAeQUgyCxJDovBHP8MM4Vh6AFXJyU1K4bOzmzX9tNM0rrk7
kVE15g0rP6j1lI/5H77r9ykSvVlONRIwkRPLoAWXgbHfhpzTVjAIua0nBRI4/fc/JMHCwoEVzWA5
ZDlb8I9eH3L5lsxw5URhGj/q0rYnCBoDuAsp+WVGcwJYWN1n6DSbNBewgiN27wf37B0N1HcrbTr5
TpCeXRaWRrI/ARxz1FdzS4Ydj6Kh8JtArbAit63Ed9sIaa/Rk5L1VZQ5MORfH0570iqBG8O2ti51
gzjiuqFbaBpD4tATCYP8AsBSYKgPah4Z6tFMq/CVQGNZ31awRCSef2Q9DA57SxnaaHlUacT7Ja7u
pyL4jFIO6nmeJrvn/rLxi8rofuKoIW9oIQu9+uc7/0MBiRN43TIjNG5wBxkxLybrQtmum3DAQz1E
pmjuMAXN+q6Lj+DTyDEjRI6TzQ5jwrcuKm8w/MZ3X99Xo3YhA61SYraC9EzYO89skv1vg/JfYhia
BIaZon6Of2xaEflOtLj+uiAqqN/UO0s+uqHYeNDTJ3DOFD+7ua6i5JRdAuUA5X5jfSgUxZ66SjJf
YNNy+ikLdo9ffWW8116+dDr2gyqwgccsKTq/p7VbWsjoJJcac8f43C6I599bHaMDTN41Bpeg09nD
JKDxbUYHOFu3y3kYFYSoYjl+Kzv8zc3OulJ2BOgOlVnmL8n17FKvWcd/pXgkVQR4LJAlUdg4nppP
RFdIsdfFnDCNJPOUX9y9ZiT1p5iqYuIMbeZaqd+WZuXgLgOy93VPZ+svWsuMiTWqOmXUHorIxO7r
Q5Ta4dr5Kol72WAtQajhhlb77jN9kKYBCOoUhlhYlbPjFUTgGAwGy1BFfou/EEBLbLUUBaXNvnL/
wVI8DlCuMT4T6q5F6wrcowPVxL92CpQAjTFgIWayiQ+VL8uk6t0gYCVBJedXZ8GeKa26YQkY+E3v
a6aPU73KiKlFomQDjutVyrPVgWYQtOegGJCRuombja0o6DYwRyIlsY+4SmLNDbAYDeyWo1n/kdMq
fXxYtXjwpuVVXfAZPE7IuaSdi7kRkVr2Z5yzNN9uU1fA/kV/Wb/ManQ6JSkyHzG1AQSJ7XABGorl
2AdjNScI+ihGrYQ2L4ZwPGc4iuAuGNCAKkZbwVlVOYPTuOxy2mXo/Sf3g5/djXsBpxBvPqE6c8yB
UN7EIZrPdRrbzqRP5/QioADFRzdSylJU3TV4gKIKah5bJWYyTjHfMdTPU+0m3hi4c0NEd91LnaNr
srYZLh9Zqe57v+lHeTEOY2A21OqtSRHb98ImK5W/AeGW6dK4Gm/3jh7rqplJkJsLiOtu4SfidyWh
Glz+RpBF9KI8kREw4yWacYdy8aKO9H39Sd5ccHM97ECTakbAqo1+o3wLZJRxfqIkz3xvMq3fp4qQ
xTx2n266HeiylllT+G9Fo6OXThVFAZ/HFl9du5Wymo/aKBQAEiYeaF/68HUv15tmL6QuYnixBTV5
OIhC/LN9yYDFZHr+Z3EwixzM2b/3GgJpvFPRGwatrjMo3VAIpQ9r1pYIup0iWpJprIaRfb9iV+Jr
tDh47iwBg3JgYzduMnZH7izSycY+NJCUhUbK60vyo2y7a4uE6BCN6Uf0u10JceyPbe4K28RE02jC
1Y8/tSj//sAOjTgegJPLpH+HFvjw42Cypr3lAKgMIbq8J+89L2Bq5284M5bAhCLu0BSvVzjtK1yD
jfPns39awQdU5pNEJiH17bV6gCf33/Vb+vNfMa7gzKh189inQMQBeqkbFKV/G9XqoFATh4e4U/Y/
EVRKySXnBEfw4g9k220AwFyFwL++25oow9Vc0hDum2X0GalU1AB3uTi7Ry2001VozOhNDiQaAC3n
3OijA6nglnX78z8B0xNpJx/E5oysE3b25L0NyI+h3+YosSxQxUr45CypQ6wv+3vMZ2fW0iKNccLy
2MguYPOIULXAVTUk5WxJD6FEOrDcxSaDwlMWE/d806yS6j7FpuioR3I1OM0v5ttOJZeiX+6lhDze
mY4wvLH1d7WYh7Is5rmeKBUJqCcns3+o4g4TMVfeJ5afAqrwyQ5bUuolqXiw4w0/G2m+Dhd683lG
AsDio44DEZlD6kwfKccsUodltkG74ekQUGw0c32ZJz1NQ8tdFWSNMc7MH6JVi9XY7QdDZhPZrsTI
XrSKiKgkXaDqSBEPCp4+ZVIaVBmR7yVlNJg6JkVTIhZ6gjRQu/knXL8lEQBpF1be8LT2sbBW8Ryw
SdgCWPda0mdDb20Qfb5AcAQt82lu7f3i9W0YwHjLwUZ9KsBoUMpAlHTqKM8evMEddjpTrpTbM2Ta
KXHvqU280QCm7N/CW16SG84B536GjY4mIR47s7gAJroLeqOWdxP2rTvr95uyEKoBeE3NUJ0CLK7b
6/+/8arsLgPhISywG69t1pObJzCengteZN5s8oo48nCITW+e9bF5sBC/HJ2dDZcxTFPVZbTg5RE1
EvshMxvSxg/wypukyE4dwDCaGlBogCW7+sPl0tQ+j1e1UhshBla3srMYxeboz/Xd/3OfRsbKbAsM
cFXjvD95BLPilRj3axJM2M/JP+UvrSSVrMCXZe1gfHuRXF5kWvvyeBeGtB9GKnQ2mK4MnXk5ffBj
AbP+2b8jj0EpRds2fvlaSg1gqtFbu5gZjJABcF12XxdFRJEmrsojsJeAGen41+5Ah4B2eCf6ED5Y
rytaYxpl30M1L08/6Wimh2Xwx41O6DyxF4hkmYi7ajhFwILcdZdleyq5NrpOgETxzybfsyhYDb/i
o+iNUL3enyadGMr0rn6KUBHWnaZt8gUd6TYb8RclvPHsxz8Dhfzp2xdWBCMTxUMhwQJMVaqynBYy
yG7oKabA9tiVDTaLzSYsSAfa6bcsP1ZxUfohzzGI5JVIjN7QIBfpeJpjjTpoLi/FpmXkpdA1YxOs
H0s7zU5xkrxAqKOj3s6V5XpS/K2ZAGAX4FNI0Sr7FDoscfuDxRpQhh1mptE97zAkSSNearR+XmwP
NaZLvCgowITWG54OceATGt6LPIMNuLaFJc3lAbdEw01VsEps/IbX/1GEqL8Pyx09L46sgLFMG80u
T5IfxXywAY3W6aHqJF6AapOf4rqehfd3uKOMzQC63twUpDftPJA1ZfPMMoWymE3e1URwtxaJtrgH
wMNTH75jktaOpyQQ+EtcKXD/OACA3W78OMfD9oCWgPx6jX8Q/6JOEuDW2KUdL7zFyUzyXbuhkZ5I
4slOSLL8cHayU9M9gcLU2SzFjDuMQzJ9L7zOmW27e9jICKNFMviDf3TBOjy5bSGAkTFwq3G+43To
cNqQ8nH0xhXhNbln7DuuBDE7Da60EKHao2Q+pgVMYcRMA4PYC20+OqYEYPgGTMp+MaVPfPBG7lay
mLu6uhB4i5VAJRca0sug4oDRSFIxDscqaFw/8Xyy9ltfYbWzs/ZSfPGwPlS36aT5C7ao4XXELfY5
MAaZ8BDdMGdeo64L7qmNRGzkJiyRgUto0d7HGO4DBnx3INWmGHsp4HsRhGLmaXuiM7ELSl8s5K7Q
z7kDbZDIuRTE5M9EQ3PSFME0sl0cQ0Q9vQzgXsisSBN4dsdasSzEJc1y9HN1a459kSvv69Z/Wsqt
sX80FWOFggY3JlEp/CmVoKuNAtUwa7EwB18owWGsr+UioBNTKvYkkviy+JorusvYcmPenuepRHwb
qoqLX3EWYKXtV8AT3PfAsBsoPHv9cLbxf44x2SoZNycbjvu7jZuC5YR7hVG2AEw2Ljdk5juAK2/r
JmP3VOGiOYpnzBck2lBph+fCkRBz+HfpMrNys43ssYYJIJ4lu+x8X2ZJJk+SYZ3ynbMbmDa5Z1fO
zlu1MymBMLAzPaydj7mKZgzso2+GdGQff0r8prCgisel9j6lo9Vid72nR4/gMBLzun99WCVrIQSA
zlo5M62ExU+p7t0ssFoBnpolRcVP8b2LvVows0s7HN67+bVL4l09NYAveJ0WU+ynyJHKFcJlCfWO
N32shWjzDdOGF35uvRy/uPkXXz3RKGCarf3kWCZ2SOwu4fTZrySF4jcsYO/uAgVWEjDXhLSLdwN8
JgjM8SmRZRezY+yfRF0oSG+gGZr/gS/+wnETHz0StVaI5JtkrTp+7C1SAsC67Tj/HkRfGoy6iTHL
HzYQD4gedp3b784AQy03fGsL/mbb36bhZwVsA2iH+7+GO57RD8FTncCmg+004GiwA21mNs9YfDdE
zVRSCLwHsEKqDGta283LIldC39GqTZxLbx4yj7iYIyltcPdjEyI5mLlRz8D6VmwUi/rQsBCCFgx7
sKclylxsF3wGldrWkDHYTbSLOpBxPGz0Qmau4B5eYtIPauloamtsuL7vdSRAhF8WtJgaqAtycDBD
8d0OKO43M5yteRe+eR7uY1INTyZq1u2fIJTI25mWRdAGaBkjWUfMJFmEsRtpAKYEh1V0gViG8zcd
hAvEa/IRG3stqH/sIOBAgkk3JB21ZY+SRbEJYVhUOHcGZAXxTSA4dHKxCb70dycLoG72D0GHzvDa
knMuphH5suZWhETTqR7pDUQpka54vueHIm2zPo4xr71R+kJfhKegybkdUe5m7LunQmH3itBcoRHY
AAqoWr6hZje8WHXfWrYX9Gt/kHF36l1T2L+9wgWCGy7XlscH3PVAv8MgtCdGvd+OioTwrQEq4Q/q
iccqE/Gy+UazzHXQ7HK/8WahXE9+it22p5lGsbu9B87ra63C79UXy7F+OszeDNbUze2g0o9oVnxV
pyJgzsxRAYTKQma08sUEuMmYVzeCLC3/p/3ZTKO1yXvODwmnTNFqJcasq4HXyR8tOLhkGWtsIgpc
P3Eb2ppOwhqLeygTGttxrlzU1hm9zmJ69IpQQtdimVdrXxOTBdcrNdNKAVIbEnUqgQWPFEKtY9BB
7+fqkRXNEGwLfI5PowqRJoNkWQ042Lj1qb3LTB0zE4B9oDSOmfbVf9vMvvRjLIKTJVkcVd1Rjlkb
VzNhEreyOpokWcarszRthIRn5HHgNmdtNjjYJOU/6dl53hHGPZ7Am3ikTM12fDyM262LJnksH3We
ZzAku7k6bEb4nLz/Q4MDEP9+q28slzKjgj3ONc1dQ74O5QjUAQKGGT8AF17B431XSjBvUgi1JBcZ
6LCtON/mRNRX7IATMmbx0L2Zml0jvlm1Qy9dDHMVCbvwFh+7kLAw9UF+E7Kod4sI+9OHOL5LN5d0
NhrsOXqQS88vnDCO7g5jkNrSHbNLaoI1NrrkNvc3dPAQ6PzHqpF2s/IwUN2DDs2Ea9gJqMobYSir
hq1vvtwCwRYzp7Gj1/A93AXjOIdJBhR7l5hBvWzMyOrYp/eAiTK+Q96WVW5Q1V59LZTJQnGXjVke
xmwJIPEJhsbsHywses5HtYvSTxT0wJxxozs8wRodYVJVmRbe+dpKA/bQcTv5FSVU7IKshKeY1kqx
wh94J77aYKFgxuz+M3XI5rKOl2EKTtJ4z9LlUlO2YVb5M3QN9/8uGxsLtsTxieVOXxZLlbY5MJMi
k3XJdiS8ZUUnJzOElVVnhMU3/KCKsUN6i1T2Kjx3VIbhziBnTn37bTOz1ABT+EVYw8g1SS2CQMIX
sJblq6cB6zzy75nrf2sMhM9Ja5qotcQQ4jEILLyZVBWfZee3ktdWvajXAj7z6CN9OU8eZhRo5o0m
XydNaMjjfVFDhuaSwtjcgCG4MXVrntgd1LK3YKPUsClqhmtP9+lS5OzyfhpR0PoeH7g5WWNhSDIb
Fssdruu0CfuS7hJP48rGxChxRtOjPAt9eEDrKyihe37AC66y8B5gfkD/3FZHdEsoMOGNKXT4GJ+c
X6T7B4it89YBNTVxukzp2v8Q7SrdDwSlLYZ/jnZ4nHJoCE5ZfTZLtSjCrf8NYI4HhDyS5bfQcLQB
yGCXLvSIQ75+jk5SpZ7MteQX1vSXu60oZ95HVKuexzJZpjl7q2U0P3ARDTxC7Q1ADwOpZTdmdiRP
9hkd7YxCp6DPN1OKSoGaJgextRsb4lU5G/LH5/1kZxmTopoApi/9ZzUzWsG/WNggwxCXG/HxcVIW
gXwlxknxdKM39CIMBiGftWjAic03oWYN/ObwS5cXdHOLWucJfNsNb342r89vF91zROkbJLllovxL
RhNfwSv+U1yK8fSO5DEcUjHjDrLvLlrjJ6728D8ZUEkrGIyr3+0IlhCqNU61ypPbhnjlbxMbZGd+
TLGv+Cz9jTm+qcTzt68SWBvvcKTGYq0oRu4eHDK+WGjDmDmd6j739ZanhsIoDlZfjSF9LUf6Wtru
XyELJWswPHD9tYJJtoh3ISZou9W2CVwA0nvSjyJ/8wx6F9ONL6LBzRYu3rjcvKP6+pDqvLoBOa9y
bEwWXw7ErSOOPpmjPFi0lHKQwthU+HbQ+brohQ82MFQbds/ysZPL2S5Oy8H5G7GsRkf2iu68E4AY
mnq3CHyW19Mzb3PwTuVidxSc2HHr69JkLi0QWqiUrmmJTUSqOklKR5nYfgcbnitSTPLp886aaLIq
isls0SoHH0a5nszd/i82LFJ658aqXI3ifQj6RRPojiKD6y+hWo7RRZirbr2G7CzliPcqheH5Uygp
xgvt6m5CqD8HkMi7o1cPX0OTce/4E4fQWe97ruG3Z2Rtw6UpmUWunyl7Rx4HMflLZm1FvruP+gMa
mZf5HBmdgh7yLtHsVhnF7vgl/00643rGhmAknfimpjbRwbayPoJgERaZt2gnWgcsCWnExf77ztHv
znSzCcGHdzUkZizwwuCWLSz12TLy3z/pItm0VdtrJC7b/dLOJC991QaXhBbK19BumJHMl4sdrHDf
6GnsE1slMsbxVK+iy2bCHgiK3WWE8i8vVcfeLvRm3eTeG/AOXVVfmqs1axlmht+BkLH2M5/gNv+1
0b3C1nSROHl6cYDyJpFM9zPe8MngxLNqxf9HpQFGfwHkl/UoquL9jppEJAbJRK8PijJ6slWD3Pq/
scu6Kv3jxVZ/DCfwV25PVlyLejrkWgy4+rVGq/2i7u1cDpoUqb0gXQZiSsIrtEHqdJaeIH34VT/I
QLVqqI3by7xBSH56AFKhhxzYmztaqqhev5fXMnd9VurKAo6DRw78qE+v+KUj4tqG+QqUMsEaDt2m
GH1jywPzCLjOsfhuTmy+cyKx3Kv+qfqiXfNuOVGMjNrWNFyhjvNDfUwD2bldugcjWQ7isBvH29r5
x6/6bkFBb+XYOuxhnAJ5Mi50ZiW7ZHuiJT6gxgIAktAOuIDZx+dF8PviiTWr2GvvbEfZP6Ovy7H5
g0DZTxKxCX+V88gGD8+UWW1cBELnTDsy3+ZCb22ZeLqdKI7GKwuVmUUDFkFRXnC8PQL+0aWjJfDe
/IdGMdj1o31f3Edx69nSclQOMN7IlKGZLq8Rik0PR4ixFDMrF9nMCAspcselUjyC0T8WXd+1wBcI
yPnaSprfaB6/58sZvNW4N+s6q9lYJPbj9cHg3PAMoZkOQrYxGQWD+Ri9Hn4R5jZ5S1J6zBLx5Nak
4ROa9heBi5V8zr+xAqNA+vEdBI+HrDd9EmwH13xURYFvCdODq2z1WHyRpUNFrJgdIKswRy1BXbzj
coRmuV+UMWEdkxpTUjjP6Kj2bAMHCyT+O+3kFsStWfFQu6/NijNIx8R1nNp/UsHbSJTmIQEOttWy
f3HMZW7G6JqSAzs1pxvj/nEb8owzZoX13vb4OEvrS2SvagVgD0APvmnr26f+tPA43t5e3/AazBZZ
W0jCSJQgXiErojrDCbYW9ezP4vlSEVjTZfErYkJOm0ODowBo2tZ2lG8/82pHW3dVqL7iBtD/YM04
alqnMXWZ48ZZMCrOiscB1kX8Vg2sJjJCujPGnWOim03CERUlgKtsCdxSyG2tX0k134qhbZ36xwqX
kBMKSdoNYsvMX5cekUidtxaJVxGFM9WoUwKT/0uu+C7tD86Ao0vNKr+HX9JiQQYmVikBVNDMEwSK
F10jBs/rrHYCCPoul9K2fi2bf3kHkmIp/48caEJe4DkRA3MmLKwopugJ3wJcRLiiWwxxXPWIPSvo
BPe6RjdPTpwuDY0oMSZJxmwav+n/hueFGdWN77r01YzoUOyhFHFHfyipcoy6J3a+srf3ndcPkBKf
0skNCzdOeEL+dQtW9/CEo5nUblI9lSXNqQRQ8kgyh0/3SOiQ+tnYMviDCCsXsPrfiNn7TYjt/yMK
G1TqLc1r6nKAIvnnltiFsN+Gj/iLqtOX0tKXvFTi5YvmioH7Ka4YQVAhlWa3mXPcGW/l6sn9KOTD
LoMkgBRxHXHu0yHIEY2eauBTF+DxUMUK9IqsRQ1ppj68MYEGAIQJXsAxuH2gQDHh1GOu5L9CCpeH
vEmgPEoZvxkSqlTo6D+DBboIzLM92XVU+6zQtADyyPlu1YSTAWwClh5RA4MBM72OvivZwWiUn7Bk
Y3FZWbTeIubbMaKE4uTQgCuix2KyyExhiUw9GPFLibI3eR731VwA2l55HfTeF+/ZvYvvhMCrJ6HM
MTyKhUDpPVUlVzqC5+VUe8rUaAKQWfWABk4FDGGlaf382z2qGU8y3p9Sz/PQiq3UlhCwagXZ/yTG
4xq/cG8K3v4k8eBYVi1HM9Gw3TXHmr+Wp2q8U0wM3YlhTayLRJB/5femQA+A5hpY1A6FZG/64/r1
LGFbNvf8f3is2ucNt4ONGwGO6EwrfWYe0W3e5OkP4Sg/TsIBmb5aUz+U4FZuku/+rHbPhIQFhvZ8
e2Uq2avxyuiooEV+R0OdYTMqHA6AJdkRESm/xMfwC/XvNH2LtwHdRIg9g7YiagSBvz21UCRaHnmL
lKqFx0RwqQ4/rPc8limmVVohEbm/7iuMdNXpDQ+Xh0YEwf8sxONNVAh8QHjGwNCK7nesK5bWRDRP
qj4UhGmFpMt5HbUZQWGNHdrohmT3294qSvjpJfrahYgcta0Mmx+/Kjz914TZRaNCu2DC8WIkVeQW
OzMJQU1/8bANn3pi4Nry983IhW4jBB/cuBqPthOeqfr+I+R3HWiCJCZ1eVhmuqMHg57zC/zfXtKg
RrN89WCJpWqeEACh12xHouXcR7JVcW74HtSsyqX+5RLTSHOXWLf8Xrijyhp+AiT7thDJCjzFYsYd
pHTnFfmTMyb8yMjVYx+t+Eaxbuakilp6wZI7hPXG96lZ4bf35now5o6dsLisn8OxOcmWM04mn/m0
GtFrWZNhKWTMzPkiwg6qL371vGC92Tp5XB12QM05jh0ph6egXkwkQgZeGbC0Nd4SXL/L7txN77r3
tcyvGHF2uYWFNaVAm0EOS0Ys/jxsL+nR6e7L+bgrSyto+nkWPG5QAsy1fR8WpGKyYDFlCBCmQS0J
k/7E+YBkyplSZzTaxYb6fzQVctYygnmgDFqNFcs7aah6bkmTzkeJiOWvDc1ORTDzl/JS6PqvfQYb
6ehPJOKnfJGcZlQGivXLJxc8oGEwEuen3CQ/lzQtMYMSsalm8PjS1bKtZd2u3SZnY+B8ArQZCfCT
ukC6pxaco0vrKoejOrBvoBySvfnBquy+8GlUuqthae/mU3C659H8pp0gO6ACenGSL5r34MN067lR
MTAJZkvsVcyTXPJBgVG9jbwrxxbxD67qdrYqfY5gzTuRW8Y8kRU4MJoPdM/TrocKuqRlcnpLI2Ci
OJkRYMiaEzZoYKaOVMnua5etsVAg1nLvvdbnvcMszxhKn1etGfcktkIHeMW7J7d6YEJrakPjwKJD
pOpvPnJPp1UH++qNb2UMD/Sa455eyMuZdDRa3bdKcMrWqvtyuBl1/ug2StOy61Ah40/v9/91cUIT
1sFiswQb8kT57IgRxDjKzsSdSiNjZz+MftZpXp0j6/kmkUy5ocpey+Nchbwnfsm6fEvN/I8yyH1j
6JZZPMGTSwxSlyOzMMMjH5fqF3cEQE9wnFlCnRfELTWYdRaWAiHBHwvO1jR3TRNgpWuVRGlYTmQ2
I6gs55UZEWQ4dEqQWq5MTeK5ESW7P8iKF8T2myA8+6ktTX2ILUJYXUDwYtIzWAnz1K5UaMOQx+/+
dcLboWaqg9lxG5fet/r7Svu+2BkGL6uL6X+JyPiK4a7eU6GsrsyCO03Iye7wSuJZBnhsDXQa/fLq
LJAsvfqRr12Dw2JZkUbOY/zg9u+FhkrcR4TjHyBjbAcYvkUZCER6Yn7CDu9GiCFg5vUMW0KdvqqE
XgyO36lcnty2IcnIIvMDEkUpk5HpcsdCdpgHnh/DH0Q8zDa012Aex717HQ5eYT5nhP5+azSPGhUS
fBzKmS5JE9VEPoHConQJzfdOJ+aVciP1o3n22bi1Huyl92ad1HSqYhFZiJM5a8HPvcvuWHW1Aqb5
qTFeYqe7rvXy6Sx6eAvGoP80gY+65uDoja+fx8AQAChG4j7xEKrDzas5vY62H8OCHE168VdSKZAq
VpX/HrH108d39TZqrtxN//LN869xjLbbf7aWb7DmP+pGfHNRr43h4B4Si/fAyveX05e5sqAb6kZK
xFqQhZspOSX0/F2vZZqz2/6BngEqSqnMX7EO7rqf3UR+PPeFq2wOHX11i1vcPCRaKU0lm1wpDu5m
AehLMDTvyvxKJd3b4NwAINWIXJsv1XiofZNZ5pHBWfuuqLkc/nCUGAZzaBz65bHoGr2c/CtHhQf/
5Nsx5uyd8KLzqTqwFrV0lYHv8bl6yWwrnvVQwfpa1XNqGjdW4iDtDXywZ284PH79m+1DETQKLsrv
l1FAAUfa7CaIruC6kjrNg3xqWtc9rRqn0S0KArEDcb5+7WQQanzhgmSTYIiOfSqGPvk4RfbNsW/t
JxLkLltBbX8KsCgCp3rtDTiZ+jpjrCVEa+/BYk4xx3EQ/8F3L/c890NEX3EAWUawlXkZlJB+7/MG
2uc2UfpIs4hLbHZjR4cOrSIUJW+4mkU5RrYEhNKO1nHvb86H9nISvjfXL57DkL8BljJxR2mT45G/
zcu/+SkeyeGs32x5sBM4wto62gUezfrSKdxq6fh+al7QgzG8KUCIPeQrNqRucnHVik6f9W6ubXf8
gt1iuyrupc/7Uuucjdp7UpzRx2abacJ4aWV4ZzJRU6vwwJdG8uX09zRrGTGxKBmjrBfLcjXXxlrz
V7TWrqnIOFW4Fte50X3+6Z0vAda8QEzj+kHqWJnWkmS1v2HFN1S2U7r1MTDBKxWn8XJt/HDjcG5V
MyNjjKctVjUSnTsZfqZm2PklRd6m0CfIERw9wr+qjjilxXOrxtbpjtRNLCCUS/g2Buwv8rfsd20K
xAvN5i/YLfbhltySsYYAcVCp8X8idhuNrKwBgZzGBkMyyJXiIYkmKqV9qbRn9X2Pv9iW2kAfLloD
mdPjps6IJU2HynF7h4i5ls64flzhIH4n76Y7/TAyUNTOFXm9o18RZgOnmUQZWlBQINkn1oASwaOL
ZZYb14z3/oTAAUTW3f3gHojAFYa3aMYXZ5rH31p/yrKUhhyvDTc/CxXaV7h8cP/7MTRaC0IGGjNY
G56B/QF6B8MAFvvWAs1zlEgiDnBq5I2RwKcu2Ym4d/H3d7UTn8+LiCSoNTcUKQcCUpcJSJjXtqvz
tifYqprZRyjqi1nhdvett7MiK7fq2yBamRPT4WPMJ4L/iwIXxB50+GgT0tXVDsIotrQ4+LMwBEeg
ti/ZFh2tvU4Sc/SWATcrC4nES7uRJBBiUft7DZPpkPn6NRCTmYpFJGOQaNRXaH81Gofmuwtc8o2N
8bW7AlS6eiJM+DB9h1pWFwbQ6cOPpdPAIVtPQYqqjbYPt2KDSXeuUnKt5Fpe7UmQe855UxK/xeOQ
dlFJVDq9MWC1LrxDvYi9+yl9Wn/w/qx5sJTM/8MGJ4Ee4K/UViqwd6MiUd6pat59nn96R42eZBTU
cESjoM+nhZVtX/2PRiWdz3+U+x0biZGthEiQRI8AtD0LePojy5Gs9NyuiIbPTJtIRdisJBznz29o
Lx9oc9kS426AUkZ5IXp1yjfZm0tBIRPk5Hyog3tExAjauSX3pHGRRJH43+6Q1NAGLrAAL3TGfBXZ
hRI/8+rTnSFvBQexyIh3YYsZSuD9zyoQaSE+khYJjabvGesXr06YtpqWKtbnSet5vL1MuXq9hEM9
xPTtHd7CSRmR6iyoVaqTTXPRcfLPgiWlDGjhAkK+c6SUDnle8g8WAoTdKo/bR0EkT6T2mDIPoe8W
lMsGl03nOMtQHh0exQY1Sjkth/6nfNS3dw0fW59zgM1wdYkt5qToz7yZfMXh4rw1SHZLUauHMmPf
2A+fzHd5yNDVM12FdJetfR+7XMrn0L0nImiptVPSQHkFGcwAw141B5T7mk6BhxviQk4lnDFsBi94
vXCmZxEV5jC6U1UhsQQsU0MKwHsVsWMvtFe8EghXJL8vC8MnP9BYCxObFI4YO+fk8dY4rjl7SLim
j8H0vqh9GxJ/AlFOwxal9EBKu/DccwDkOG5UZXyRH8vogK+NDO4IGg5VuR/kQw2UKXVcUEcEw2n8
td+vgh0+3cVgoQ8YVmNYkL+10BgjFxn8FdWqy4mT23mSu/AOsX19RsVPSwhp0sWAIaGZkjaXVErj
YpNPOwbbgx/VCOx9oyqKvkcOcADf36R545E3IIPx0AQhSTk/ATsXNIoYr6r2rpywTAF+O88cfQ/L
ii5RMoDN+r8rFJZGGAHEDBzNzHgDID2Sj0vbrXv11JbDgzByhtAyENPf+j5+fdmy777kF6RU/mXf
IdetGzJmofzcInhx1up7kKB5SICzcr4s2v20hG7Wgb6MuDN/W8tdTqriAU/2UxY8ZbguqIiS3e7v
7EzMsW2/my4EbOOJeTSsh3suDdXbQdTxTNaYtJ/TuMaDuE2vR9PvboCpXskGuhgW3ts6ft8sm69u
251rsvp48pGG/c0x+DorQlELEwU3UoiCemGrmXhPH46TYsW8/FE9CfRCX+cIVpzg0WR8OKrgkLI4
jc4aWRFVsClWG+70A7SE4rEX3KRoHburVd+lLPsDU/OWqsaR3QbBGUAzYQiC3kRWpezDhelSYyDM
Z2p6c4rrMeNIVsQLAlFkO4LyeED3v3iDxHwSvWnpxLntYifOwJ3VzRtjJDJxsO5vrz1OYxQdg2Ke
NlC85kR6ADo/PyUpBvmg9zRoHBEYAvuWpEyNtJ9J6IXJJxTOovqXJ3uP/75GNm1Rrh8Jmmn4w3+x
eHVnpRxJ5A6V/loMbKdrmbyGpO5YTv69RMLbcIzP6ZV7TSDvTZGvB63IDsooF74sbFsoMEx9jVe8
HZfWL7dSkzQkYURcLILk1kIeHvaPt8NsT+NA3/bSgeb+parz5wPrjynDqNmIEu4ax6tr6LU1TRJQ
PGMwtBo0sIzZYSNixi8i7mp3TK2uBrjkPhczYnze+5izZt9KuoyJqcCMDtx/iSq7Fs83vt3C8ktg
ZMQ2dO+L2iLJgXEAZ/1n8AKcTFDx6DS+5nmQU2e76hH4LUCx8pti77sqdybDht0lZLSL5zDRct+U
xf6KQXU35X1mNmqax8ZiZ/3+xSI5qYKYUQVyWHJcp3ZDIABxL6A12ZNBbZP0ixYl+l81BKO311C9
5DdcmR3JyCjQyAF8kkCnR50+cRC6q3iCII7r60eu/qumxRT3f/GUdsv0kofjpMx+krHRmc6y0D8Q
SZMwvWnTFLOd65bey8OvxhUXEMysA+i9n7WsSJXfcVXD1uhgfDgVo4of9FbgIBpr17NizR/3WIGs
wZ66JeQzRtU1YGTcUf9aZnMGnwFeURerTQLz55T7N7hVOEnaLitm3/hVC6AyJwoPx2ACjcjMFsrP
xgDfMPTRGe6VCqxEsEZylhk4TSBZuKYA6k8ygTu5Sa0UZCH1otV5oD+FdowSfiu218JSTjcvUnp+
J5Il78Y0z7pqjKgByPHsXxJA+oqViTmGmXM+kzPUMmxIIJO70dMKrxEDQ3MWzgTTO388IBwgaKxZ
BsbDDixidBboG3Yhks+PitnqfNBYIQPRDWc1dXkXJc/vZ+aBXZyHilXjvw5IYnyXUePtb/fxeRc+
RWI1992lUCFDd4rkXFYySFFFUubNeR22C/5oDCy7B0gsw84ndPlqvHircQ8tXt9NuF1NG+Me1rZz
6Sq9mp2/VdvMiIAT5PG8coHKu9UoK30OIXVkBoXgGYemDgNekJYeqLzOVxW7UsJkAj0o2uLaZmJJ
iD3yS+9orxCrnuXUSelAW9U2qmml/WXwvjAfwD2DGrzdBcBLgG6S29MuVtNOzd62eH2aq05JmSCJ
Gpi9Blhq+Eu1WHShp5MNNHXwXZH2SqBkZ8ba1f6AOoAVSA+5ZvtZjlYrAKcq0Nek8vjnDSAdL32+
ELtXhqcB/HI8NmBBU9JKU2OP9tDlOWwzNeT4wLfep83UH/upChnq8aRc/fBF19C+Z10hVUE8WLK8
MHEyaZb0kYKz7fczkEoklIIfhi9q236qPM6WjD69sw3322/H1t69eGIB2drkSMDocNEumRb+b35O
atKPzydJImsJ+QHMsBFmBCSwmhvM4TuCWc/ZLrUacBk4OIkl1pDBR1WasPiaA3Jw7TowBfdLinZk
AlQCHfxaZYBmDBxS0JGaGxk3N5K3f5DGcbkvMQ0Ss4/EFQzxUY8g/269fv72k8RvUFd/yYaQDqeO
Tmi1GDHxiwTg9cfOcJr5+WSl+qfWq03ShMsFLls2YkRc9q3psacmi0N5L//UOrbNgPPAvBIg/HcA
+TaMQbLjciF/w009oykjfePQRrN0youAtLS7HWScwPLOwQcVZiustFF+lInbjE8lPeQIeipHRqIH
myVWS9wtXmJJqNzoQUZUSJwImg0SC0k5mCEaKSMC/zEy9phr76KPIzNKdwqh5NpguXNLtXfku1NK
obSZ9w0HscWwYpqIO3Vg2qQekqYTVaBigbaC4YAIEgqE+8DRW2c3A3tkTSp/BDeUaIAckjL1qYlK
TZkmAQUt7/JJcZ9smXxuYcWTwPyqSbp06KewKFaHqb3+4ddSODCmSCqpTrKY+13ww1DNaYNvl6qm
XIjOh5+f81sIFuTuJIw9ztiUAWdpu2scIkzMy8F7Ob7r8Qc+NVARGvwC3itItqBY/hwJTp7Prs23
LtPFgLVD0C5NT1Tm8k0a9Bc2TmrO8EtRoIbTk8qC3auL0YnHI8OqVuOaUQyEVnYnee3skBQU+m6U
hScGPzP9upqGWKlJKqsvhqWTIvaef+VZ0tPxjOSSaszdCdBY+J349PIXPKwCMiygsIx3x+Dy/BES
hZPStVCTWVeVrJx7fgrS7/nID44mRA7IAxB9tR5fAwZTy+HfqEK1nY6VfnI7/HVdHOPur4sWJViE
MRD/q2SrPODNXgf45gggYpS6bsW26paVI+6au2wxHc6uO7bvfh1CNty9ND5nZnTvdlQXFEXMBzmJ
wi05YWWvbX6mfEi9YwYie05FMsZ6Y10DdXmlqzHl07dShh6RbbQUk7q/JxcEwinIbr0kILh0J+hs
YP/8j1wGcwoSlKbTNZlUbtaoyN+sqrSpjzFimppUcjbJfbJJYi2OiOGniq4uB4Aj0DfYgEtQ4Dlj
usQXJ/rZM7V4UlL53MqNHjTs7dGHXBWxLZOT9XQxkpAyhgoiw1xGwVlxSK0FjnjR/fPN3tfJNYkn
zJm7mNN+69YO3/mYY5UZm7EA9v6vsoIClErqBld2/crUeQRoCLhep5jUGm/wnXpg/JHbiQCjgQjV
rdP7gJ8LYiWTwxbaWbLttp4UOOaJEu9EhGMHxBp41SeEncel0OIICblzm8bYzXufPWmud5UG8X6O
7ByhjH1mBdtX2xxxoYFSYVyNTcfM+rk4wCoqjs7KU/3iGgzqS/p7N20p6+XCFgzd/caaa4YLnldF
TR52N1XErwLUfPJ0Mbkr4HqoooXutWZfZmOWcnPsIKEZbQh6LYUKpwco60oj3PXgGZMpirLZOB/A
Waj5xN1AM8O9H23Pqp+c9RnIJ2fqZksnXkw4lpIn5xWo3W/nWFN66NYywam9jkfZpE1A2vZzzZ7T
U6KbbThIhUPT5cwQWhG6P627nIhJBnokD/GbhJfm0IpmUdUR/OA4fN2SOksEs0YLN5WP+Dl96/9I
3T5lA9dXKLBjyLLgJemhhqoke4ZTZq8v6Wki+Q1wrCWDvbv2520eMimyJODJF5EHwq/2XmQVj5FC
MxdP3BvNVAsrMpbmC9PzCU9rcDl76fZN1EXuEUj+OoMpHyV9q/dDv6mDyU21Ho1p19g4rOQuBe52
suVoj2muGyy75ZtqWIra2hmr3zrACOxoHYP/N9GrQ4EbxaKq7iyp+ep/E70yrcEJHKXaYtl/Uq7n
oF453CYo/2L24G9Bs/DZbwSWm7vg47hwsLiYvjWpWX2MIny9UtQceLL8/fA5na411a138irv8iaC
S8JDE71XJGFOpBc7AfAh0P3XJmOYEYeda5OEcJ7jEH5OCo/JxG4PEHF3+GKtuwGGiqHltKCOM5Ml
7iX1hxZAQ6UG9XM0jFnOomFHjy8bm/pcZJ6JOhTymO3EIyBEJG2B36cz1SjCZiOMoQcTkzoFB8YH
3iKG3Mlul16vjkuhAa96XgxDuamW1DJvHvywVnBtUZ+JoqWzAQtuz1Qp6yN+pYiriaZ5pIY8CYxX
8uMydkTa1Ic59PVPIOJ6Ue0/sgbiVbCLE7D6KnM7OmXeey5EgVw9nWkRBV1tHJX6/+obE9QXOGQ6
zuNFWZVyp/TOWiCMCEIlbhXop/sZvXCJllzobnEtrFfNx2wR58Ejaxv5/tZz4LzQ8iCzCz2gmoi/
EA2hj4GAAmZecRJNDsqjxVbYDMLpH6GYAwjmU50RCv8fG2d7OfL3ifFJx/sMBjTFHhXRvC+lqRmP
W1sc6V29bFE2hYzYMFLOGv0yRQsdpT0qQMbIADw/koUpZm8W/syIaci8PBJGWVLZY/NkufBcsXHU
solapWlCo4P0DH32KOAaROuJxoGoZMzmSKWQkQEguPUjGObVGlD8IG3FzVG6i4lne9vhFDNCnigh
WYjZ0pL2lwCztW0Bj/RMqDok0Dx/3GQIKd2t8DARGxQleaQ/sT1i+9OMVxucB2WKNzCCG8M412PS
f12MtbSLkw4d9UCtR1XfvL08Ekku3k018BJYi6NWHLBZi/Am/Q57cN3KimehKc7WR7AvvI/4FFqZ
9yfP41geD4jd7i8tLLBXPGm+F9a1f5GcM3VpJPDlcPF2SMsxI6ErIqC+shKyBFr6l0d0psN4l5ah
MnUC03gJkQuUb9Y1indzYNWbZ2m7h1DEyVuTCPwpbrMaZXFHXUn8j4d4lXOb9BolAH6YAbJ2G82L
f7jf2q49BXqvevPlz2cq4yuFFNEhuaYPX26XbfjU9Rl+txE7VxiWBkdG6PAHMHQpE26uWE7gYwNH
i1Ql0IHBYfI85HAoI16UwPha3IKh1qxkzP7Ju57QrZs8z7At7SKoOJ4qhUGYfGx3TNrOlLNfvShm
Wn0egA39b4er2iHD+w5bNz7Pr9nq1R4QjhmGhZN6wodagEYt0VJV+AUsGINReWN6ANOWXYfPHCGk
eHhlKGlJTIWQEvyOWAenggA5rtDNMI6M5CRX+FD55fDflKLd6DCz+W8HkjZLm5U6RDouG+K9Sa+D
BjWWnVyRXgm9GNUXdtC6HwJ/81d0SljQZHP1urKi+jpFvD5R2kmRwK+ynyD0s63CRTVvarRJ0B8V
t8xOvJaJnfu0Sd7UBFtMGNoVl6cfv7lrDSpsTSWikGJ078Iin30uD8J7LAsJG9Br1/+mOYqkxT05
xtcn86Y90hYIH7J0pQGMDQrA2HziHCqCIq9igCRfIAFvJNEDUQIf5kwdFjn+oPsnRK7hMjfDWbLV
tjWxMiS8B+FY2C79qZqsE/l0ZczOi4oG0RQxbzw7aA27mbjdV6yFRgE/gEm/D4kJOhAH7p7wBYFJ
Li8yroCXwqg1kpjNCmXI2M5fkl1HjKipqrVwvyY/GQY8qN2JUHmQ1nRkaAZYvZq+cHnx2egwfOm8
STo4h475lpa+mRLFySqXGfSDbuJh2hJeh0In16jrOgBRAMErq3zzy5xiIoLZiGMhadRbpmf3OOWA
Vb16e7kur4rO6+TExegwbbetTmhWCa4i1pwn6Qsmgiqc/VVi1JIQxFRIzQJCInMO05Xm5ZNPOqcB
k9a3ykRuG/A/oE1hYmUDrxxn/iJ0tRlrkYgi1sVp9PfXZAHwjoCvj4OlXu0ColGcj16O3OncFtDn
w/DljpshaDJ7tH0ThO2QrR4a2b/NmRp4Mrf8+DaPxsj3UOVlZG1nwpMOb4bOH2U6lYyS1Pfc9nex
BaC1qVZFcazimKEB9FnVKLM+txYH8sAV7bTcEMsYQSCd03DdrDyMG5qxZEcedkLGpyebRymsIZFc
BCEuixL4CHLkKhTVWbEFm+y1N6jKnHwuvKI13edNsxghmIG1nDeP1FKejfxG2OvpWt7SMU0VXcWD
NPH/E2h1HhsxO8WqiDmHIizQqHO1Q7qmWcdX1OurnfvebfQId0PREBYV/h4FaOIrojbsneEu0UUJ
bInnBNk7XCO1UuFqGnV3XCdTuGgqMyXBUUrRdOkOjTX08TgzFPFgsP2X94Ob79jXgN11Oba6/vTK
LWw7xSjXSAqmwqWGT5lIhmBhRMKsWctwhgD+1ksRzWwMuCqBKMbLyClQjqbLVjcSWz8nxo8RgEMl
CbUVDMecFRlDeh1VVR1KiTptZG4BWnoLj9P0VZTfI29BLSUExGSfbJC8anVUUW9h3TVi9nEJz07A
qPw/7rimNWoKTA/E+OEgjDNt6SSlukaVO3z1erzFFla1+mOLlJG8rYqhwd9SpOvucH+vpZ1Epo1Y
xNrM4Gh6glereR7iMvq61fQvj+19PhyiOFQ6cQcsk9VHfhXeTMjNjpkGlt7qX/n/47pKc1dGWC7A
u9Noh6NZVXj322jNFGTohFOBM1ECjT7atZchyDCQcDsxQIP/dRRD7w+L2PjMnN4iVDZfo5/GYeYI
mHeVjwXRlIEVgILb9z6rUpbPDSDMIz8a50HeOF262XfSQegxeyCc49harrTvsqrUdORY8kxUEoC1
nPVNZ7HaUHvaUsmHygWwQ6y2tLMCs8n41lDRWdIy2yO/nqKmZcDJXVewjNRXCw5UHg66paISKi0R
LsZjdERSEb5pwNoG/E3CPtvgYSt36kls9twIxdG+OqWxiWLNJ0YgtwbGx2YS/lgyrQyz7QSCKeuD
K7gKyjSpOy7BfpsuEvXaolQoymz/N07IIW9bJJu2jfVTRm/LWJ6hCIks+Ps0SOXoeGlhXfHhNYjr
a8Pu+tQB56VCkRZRXBsCl+eDuNT4HGUAnR+Xyt+473y/rOiSoXeJoMKAm5suxNz4tisVnjwkjoN4
6u16zmPGXm1uWEqz5dM+8HxpSTSxyYwGUdW4EXelmohpXfOUuP1kpWdOz+24N39kHnK5M5vU4RRf
MYKQvcl9MYXXfYML2QwzrJ02SBzhOtIyo1Drlp2ilAI3SjFB5pHTdC8l2VXz2ERBsqYxtACqQkET
5m0fOO6U0ZubWE7Monqv1dyF8jsFg54SC9k9t0qryXraXwJKF0nGQLgB19IpYmF0vJZDbcewgQOj
qhJC45bzWP6w7q/wdAimw+ZhkAr9/aeLmbyEY1DUaIKgQquVNJE5/6LFsvwmWsn6kYgWqxqPpwHc
cNqh7AV5r/datkhN6actV8zhDYwXj75imVXFToKk3lMgyysORHU0+9vfGjAl1PsC0DIL+zj5bAbO
8L33WAs6GnOAVxJ3/sQdA+2d8lU0GH8/kEMj7dzmZgf5FSeYsWY0Pzwjaarx6JcTiWzrMH8tHUpL
rIAhIHoya0cjAqsT6iqAOW1vsYOhfYY016LGZq8svQuaOsKol3nJBxdWu67F4y0yYFraPuMqL0i9
iJjmOySwWxdoWJ/ANGLy+vV3uxjjq8Xy5JWfNqobNbABwLcVwUIjfUnxTtj5NQTwqjVEVuXW7+mc
Fy3HF9C8Iv+fox5V00meKPngmRQPg8v6cWZwwt56suXOybcwttVdtlwahXNtbyYxQ3hC3xk6rYv+
3wiMPk3KeEZdP1iBwgw4X2dOw+rwOBItaowjcOnG3AqQYvWH13VCbuA0d2kGGsRnJxzN5kl9Gg1f
THSmQeT9PJDoUB+l1bpdFfzzzp1RJ1djb+jDIerQA2bvULblXyQ8YtYh2uyYZiQT4Or/h3bzMGq9
mL/MaIlEx79Pt4z6v9MDck/NQ4ERQYnGrsBvrBBnyN//vFpNsTpSRJxuR2CZZjERkj2YI7PcWWh2
o92HxqJgz3SGxfcJyOSoGwryAwZkbGd9cJycRIRYmY6M0X+M+fjnhvEcIrnR0+WnKWzHDS6Mau1O
4yN060zWIPpiRT/vOXIQgIpdSsP1Bb+YKxbkwGCJKZ7Zry4RBJxaq5qBD2rQprk1nMHyIYFdIy1j
EevEX9CuGcTjTF0F8SkS6PRgl0RTOCsnqzGSiyRDjmf61x+HWfPNjmhNLcOcOOqmwERddLsBDG8l
dCWXWGtRhREz+yYIYzNCvw8kX2YNkeW6pG5ncjgaqt4pUV15DcCAOMMf6eOUs+YIXpjTAoDNaapL
iziLvvkTYmDv+uCNuUvl86OEbqi4pEZMWqdGlJDhUzYTlJdFXYXgNyF9X2ryodrjD8pEJ/KPdNow
p+f8VHRLPLXULmEYvhuXkJpTk1EOnfqh2wRbfH3XxkK2s8stTBFD/T70aBQzKVz3RkNsSmmSBnEg
mnxZLbKL0L9k3BYPoCCY3pF6TP97vb07khUv9GQsWdis5dX/Bxec+OA6KniChD5fnU0iYlMurc64
uZL/459sd4Q8stK0n29g/qPnsTvFEilXsZgmkHzfGVWjLuCvuF/Ut/wmNKkmJCnCuzHALAyiXQEs
x94rWISu6p7HaLma45a0iQ+WobF1xtmgrpF8nmkpCcv1sXigMLE9FfeA3OvXwu3Bo6sAKUKnOF4k
0Q8o7P2xFndAOm/vYH2xPRHe5nK+zdAxC/ZjX7ctG4TJsFDlkEXKrFU9pd0S6fX4VH4SqGFV7/qj
C3DExE23im+jCjrIUIPzn4/PzYltKVn5bvEOv8+XcWUef9V8hQDgKtu34VUTKnemKN0epZEfVkjN
eXDpHefEdikdLNY11Ucy55FPBB+EjYsGi6/LmTC5gWFCOYtfxjrQ0tqoZxb3KMLxPde4MCN4X6i6
1MNWCez1f888R40J7clEknMTBVmgLOF7NkEg1zP9o7iksD3uiBs7Afj/dxcrDjAuGEswFLCszU9f
EQ7evP6gM8zgWsJ/FfWD9FeoOXHDRNirW4jZvKgJbQ/QCPvmjOlTnPjJ7ph6sh6nnpx6vCsentf0
faRkIuwDKxZlXUaOi5FLqW2S00nn1sa52Fikf7HMVhZBRmCPGwakapLL9e0+TZR+8rh7cssrPC7+
uc17UiDBtOZ1eWoQTY96Lv72fGJXQwoH7Ok+GL4TqmlBTWAb38pk8ezzJd9uus50iex7xWyIR1UD
AXaL4+Kh1zIyRW4LyErDvYqnFGllR3j110Aa8YDcQiQxQQaXktTvh5zB/WherxqH6l2P9+Q6zndT
84IXijngq/D3piwizrbsbha5Agal0XDyccU45OKWJ8dCVgbwEHJZJx5wAZiApgS1AnKOlygFtF2J
JxFJ7mAA4hZeZNPCcRFWHP+jBjLUDSX+KJ1QwTM2nu4LpPokBt7WRUKPqUd0OPPnlpQ4E162BcWc
h8LAWbbs/tyN3DYOE1vUZTgUccvzKKrodpIibBDhxMBTMTNkbE7rl4yQVvEuYhWNfx6ypwWSCnWP
Fg5LkVt8+r+i3j+RW+B0r1rZrALX5sqHpGzF4gujIQLMtzhxAPfMNmnJEOOrdXs7fxSfmlWWhKkC
8/hnXTPqwlegCH6X3OuGqsB2Bkg3+tK6PygPOPfZonheH2zWYCVqe1wOMlTbE1V0WhsuduaTuBtp
itRmxbLNeE55aQK7pdLN07NC2b/f8rsQ6i4+IqxQKG/gOkUEByx3jX95YNgCC9F3uRW2zk3v0HXy
Qq1/8f3n2pybchp8NTLhSRoD5+cB3XmqqRa1ruGBguD28yki+qXYG/lP2B6d6/ETZQ10AY0fVyIu
l1qMDKdh9+cLly4ExQoTKrkGG5/96yIKKxN55MkbwLxU7UvXPE/xnnfxbuHgmfDkv6p0UQPgccKN
w1QUWdvKQJKsPx18hJPi9huLjurJ3Ruvi07C4nNBi1m8Z3Q+x4mXtZSuUn4BwyLGB8HXZH61Pr10
ehYsT0pLAHDqCHpiW7lZlpm27Unb5Gj+y8Ygp3YiAo3wSa36hnFO2RtczIifyX0PVokfPjloXyBK
b4nu/e+6TitnO4nKpqhFnmd2wFZV8JW/BvURnCtUhoXd7QQ4gymuE8witytJvJvETKo2iqJZzehj
VbleQp0KBQ4oWME6vghqnQtgQFEzRPnWL65j0M8aFlnGQalzCQMyukh8U1vgd9wEHnwTdxKeSTCP
t6zjiiC8hze2au8HgUVHQeFXgMWl3/yRZek6ogfYslOzp+VSwJqZ867kmJO7Iuy9vRwEh5JqMOA8
0+2v11rIxfiYua/XlK7zVwEm59zb+NGxQz1kbBhlQpPxH2euHAPp/0n8AoSHgiKOVnrxyHp/Rj1E
ECDUAis/4opmfWlmQWDomcGFK2EZdC2awh0mWNuaLe9AVKL1ABut2ALKeCvYPVU44Qs3WzYDjt5H
Kz/qdIUAZo6wTq8spV8L4UNgMXr7ehq/TrfxeJcF+inwmG306ORGYgQ0yCdWMKz79W7Skun2hd06
2rhJ5Ti6vnJqD2yx5UdPAweBJk4BmzxLeFhuF5v+0x7vFseNIrpNF/ECsS7oZK6vd/5CwvDD5sZl
rhU4y4/KJ6k6cKqBdT9J9mF0L5Vgg7cy+Cc2SClxcEkHI0btQ9dM2ZZcr0gFtv77UXaM3T+J6o6U
vZ07pkGl1j7ohrprK1kULrS23BG7YKKyiPn1Z1iLx01/g0BFaN2c0hxAVTBRRaxcaxJi29cMp9wj
lGN4QCJ0yZPEYVf55fchEA9FW4be6HzUsTPPOz/srvhy5bDl60tjJBYobYJ7dHGMNQ/xlgPQFwcx
MRU2sISSbjghGfhe0sdZb3FqZbD0MHtBpUigLCZHgJznPbYlrkOc0DwyiIifPOMyzxIpEPfNUiIo
xwDMbItVsvtdifBF8Dnc5Qdaw1e0Kc4uVvP4weU4h4Q+GAfFyJAYCWZ9QD7D5fAyfyDbQJx//9m4
43Xt1W+MdRmyPwLE191cGJAtsXkIN0G9VtqP8hjmzQ7AHxqbdaRS8gveyp3UELegYMr1POkQ9Lwp
6a5zy+fqjuPR63N4Kbn2R7zHyLBpfmxRDvYqnF+mW9mqottRk3+c2m/GsZcgj5Qh48UMbUVfBSfG
Q7iJLFYce/inH1oHrU3Z+vZYxuhAcAbl8CO/+xn07YpeD9RjwiIkRVvi8rBMP4hKIoDGWeVwDE7T
OXbnse/6fx74yOjLK/ZCXmp7fwGe2eVHjk5NLPGTIRid9HnjHwLMuEJl92pDYaHCCrCCYBlW05f/
7DoJjpwUr0Ipf+5iTdC8lOJAdLXTpLtu9jsy066pqaVsYue11m8mF1noqZJCk7DGjD3R15a80Y2w
Esl8FiIdzyqRAjzOEEsoIK2UwxQuRgpWZZS9noKPgQwlq4ejbH8HayHRCGGxra4y0gaEuZekUthF
5rR98KxHLh/zEnC5l8KM48mtAg0jpu9ZnqBTXesKu2mCTBbclywgHdUo37EamlPsyD+R5Sv0nirA
/Pa8tmPGdmV6ujWJX1LMnzRli4bnks1aK6jf/Su/iZhp5FknESYZFMlDAW9+luC7T47X8/jWh4Mw
dWE7NYU9U8qfLAG/Dc8duBjb9ZgkDJOlKH3+sJG/zxVc/NlAolyo0ltUlv7LTGruDD+ISCl3DKev
lD64L+o85IE8XchL+nz6UZUBIGwBHHP+UaL2yqrHFHV0atkffyfUFunZWXScLpuo3Xs9NEwYZYnV
1FwgV5/hG7+WzBSIHasR/aI5UrXSU/hVS3z+GIw+sMu5YcQ1ycTpifpd8sQVpDZlmsKSEqXKgvCz
fZuW/Z0iVYW93/uFiCkCi+U1sH2uunkAlyh0mVzLKL4mePYkEqG6aDA3xE8aoCrDkH+RwCqUcH4p
X5RcnnQd5g/88NcjpzALG5za0Vlvx8P8aFgwtkGkElSICuoN/pEes7P6qDs2v7TnOmfx9X5Rx0gP
Hz6SKJs4XjaiXmF0HKSSHLAOo+R8U3n9hBuCw6wD2NMuDPofzedOg/zLW7Cawy8h0MzHVAQegYUA
ywJ7NX7NWB4SrjqErnfgoooBNX6av/4p24B7P7PVglm+kzE1cEgCnHMQY93ITB70mWrjcg96sYwv
ma+GeebLgmr1ZtTPs/Yc9nm7/EBGNnj9an1QoiSSZZuU7VcwL0XUzhB3h9UlZ0Pnwy1dIKeAEGd3
L500MT76sd6AFstgpizb0DK2x8q0iuOpMZqHJGC35cInvzK47zI5Rfct5rjkVDyQoqXQVVV4bVsp
wFsS1ZnZ6Ph740CzwYJ6M1g+0cbVhCUaGWpq3IonHQ6RL+yAAi0O6doAvlxrA32tt2/02KrYK67G
NDlkGyGQUtDpqXh8NWBfJZbIGYSZQhdPZbaODx7NriBRHvEsmQGcQ7QSHZeW19vHuAyb0ApokGPC
TuJmezXxqKZ+ohAhDYsJA9vLfJyp+jmEg2455YUYzOWjm5i47/c6irFi0ty4sZYs4pEqAmS6PXd4
OCy6CETOYhxNNnjqsqUSw1CIL/swBIKGrVwbfd1DC7aJSKyvGspOxT2dRsZHyMjObJiVVtJbbTQC
1UcQBdrUT2GlVN9NMzMbfI+YzpyjCkNecl32g8j0wpDtPEIlwZew2mIB4FlMmUjtwL4dao0Wepfa
UrRpnkCowv13fA48ET9V9/v+8v394d7HQbjmOD6qMfwgbzX5Ci50/RWYjNmATaMC3/WYrrcUFz2Z
KBl51Gp2KtClWguAQ1Yg7BZdF/WfsJQvignk2AIQYiPiwNFx3ZTLkGN3hJN3/+Dm34BTjmDCD/8/
GmfGgga828L6436pYCHjL56U3yXsFdg31to1Kzi+2Y9/u4ExLKIDObCSGFWctZm1Ec7vKmQVBAjb
/wROrHCGQFHuyU2HVhUXK31/7OaKq24Va2fBKAYObUILgrq3GKXBlFkloLEx/DkZ0rS6JjKnfQ0P
qrNYt017RxT20VmLqV3ftmmIFWy/k1t1Uqwlxz0wJ8XU0OnAmz/N6MmZu2MCvShGJ+krY4u0PeJm
eCk/0/j4ExwHsdFlZsbTSA77QRFVyS3zhXr+UJxsTQ8uqjbagYtc7JVvdtuuoBO0hIyBOfl5hgpr
eCzFu8g8av8DpST77rW6OoifCHqF7FG2hWL/fei1Vn6kuzDeIkXzt8djlzLOHQAIIAR5o9DBMrhR
e+xnHvkFh1q8kUaCcsnziu1DNjR6SHjLyhmYZiyRjYYK/9Tmmp9gCkTO8RNu9imWs1Uo9hp+Q7hm
w/26rB/chybiHxt639jgoptCENWOzJU2Ive7TO8mBrzaNYOtz7+6idlmXy/iykypPbo4Ry7Hd26U
6bfEz/UYTDvF+eBDlDDLRPpCMHL42rylXE2Gj6m0OK8YF/Ks1vhXSgimbAHP4HYIraeF3rfgqWFQ
8FNwGBsrVRGllQeSH7aFN3gqEoO+RrmqQ0SjzqpzVYeZrndtCUNtJeTwxvRRpLEJkBprO4Li/Qqq
E5p4LAG/AVgPxomKbYipAPAczSGKbgYvs9ck6M0cyUVkAJgG6YMDcWLJD9QlrYW7JJ9ULifIi2pG
Jusn5kIKd0brQyY5FQ0nTO8K52QE21QKmNYBpw7TcJys4Z1llDFdumsmA9/9iKzG+t8w5BQi869p
BKgGIKpSVowTkuZ16aCCxU87kuzj6GCicVPmYpGsd2M3zyhqV9uKOzFYie1SdGLiYLUWpBSl/QVA
O4MXpJy8O8VdXjxG77x4a1h4FvpJXuh3bxAKjlDERzdVf9kd3ZE7pfp8qxKaAMXijYB60cCK8OEU
LVSZup6PBbalGvqM2xoKHvdLxPt4s+vblT2wwetWzQudNILcwhV0wBVBqGq7X40fkLEyd8+YI4dA
421esUkyqklX3oIs9UWuSPpeKoXVdkSOt5IHfRgY5OSeCZD9lIvrJd1R//ndEVFVLi/x5lZM38IX
XOaWKrg3CxiXvP2PrEDeNnOvpAhhWWFhIDi8s0n4dGsHIpgtDRpvq04qv5YMe7xAZ8YT3tCpsfzN
5QwStJEI/Hf/qwFgFag89JVCXU1MxraGmzOyfNWpmUiWkB4vJKcKcFF2EN8ssH1kaYamWeBcPVqp
5RHDciLEUcjWiMu99oq9hgIKWEovCQ073d3a+6nNf3sDXSrgGd1sEoOotjuvXATHf0j44EEzZzgk
M5dKgOiYBVcHVjAgEbpkMBbEiAa7vpmjKcmDEAAOi3Z+APLap713J6hjeleyPs+NqDlBaHEyShEf
JVn36TTGLylK3O0Tmg8JnwruJEO5/+8ThyiJTVPcf5hNctgV31JfNjgDO/l9GqctD7+/gJLEy/EL
5GSiawcBqPOWadeq/PGfAYOhfb2JXK7A+6RgcQJM6zS1gb2obBEewUhcr0qUlNqhTibf3ykTTmbm
I7QttatsQqmKTcNR+wXOOLw829Sru/R/FBnobp/eq+TQjpNKr/tPsrSn3letJkyoB9DzPWH7hTOj
udm2LQR9hIZ4ZmjL6S7zX+4xMrdpjc6/P6SeiQa/buRpbrv9Co+1IVRvaVjOL0rQevpwwEO4p7G8
bbwAJNzez4umdVp9LgIARcQtIteec0MnOFZElnrNyDyETTI2SgurSy3/+2fJHWsbpZhTJIejRtWd
E7FVEgKtAt5eysxhm9wQwN9EIdCzp9qmU4huoHbcHvD0rCnSQ3M+EKJ+xvDN+a/JUTcANQprMRwO
ywZwknil86cBBAG5qeHQd1OJmHa6Voy7/7pVGAEfY9qGr6M1kOQA0Y7rZiD8//daqvP4gZY9YY82
IOA1r2cDRI/7IqFSOausEFYuedOj25Ro132XEwCnht9P5ZZFnrG4Y7DpiHjWfOnC1oUowGd/otJu
fTXzCKksnZ1Odo27OElZTc+LYT5IltdpcLOxlNCeaV7y7ZVFPkLT9XB92z8oeaq1Ak8MQV/N/1NE
OFJY4kF7ZP0LImLCKv+75bHQszfANWc8EXDtS1uuxAkjmvpxddpRbGMbI+t62BX7R1bS3qlT/Z6k
Dw5lE4qYQrq409r/zFoZfN30kku/XeJYRJ01OCY1acv1Crs6/FEVT10aSUsmxxmRo+D1RPjrv1rX
Oq033a7oBtUtA/r+Og7WKCf5oabf8h0jEGuIv5QAAwaFbHTaTXMYD9iuunTRGEtg1aUXWs/QUp8F
LaciqlJmrqo5wKb9v3SnQMm1FGUBSYb4VnrMaQGiC5oP4Ehw8omUGk+fJ5tbiWbBXYwaypTSDVNV
uHUzVxd5KZa5bah53KVs5DVfCIyrkxxK4CaPBZwdty+9j53SiOpvevfyt/UPpX9EvBPMbYFbo7VJ
000Casw08jV01vShw9z4JJ9dw9gRmu++If/jojDoYKenkD6cxn+YhlIudqswdyb3ttuYCJwxJHv6
7f+nFPhUO/9MeOJ6wY4AUepF0krDw/CgDIqLk7vC5N8cBqXAqCC2dtDtnfm+v4vKoJE3chQjTvfM
FPhSARw6sGldt87r5/Ujtw9hfdo3f6OUUOUDJO31syiVINES4Uyb3yJRLDgw/y4gEVXjZzehpaJA
lYcNHol/9vkPBmoWn6YAergx7ER/Ft2/jMiMQ0nod4i6xqptn+jlKikW6d6d0AZegrY8c3azNXWt
hcikDzNGhCwKx3QRFPrIECKmeKBgXdk1i+WqXVk7xiiKTXY1BWt9BxpvSRua0U3VotDtMI1LYLjg
uBjzDZiBQKs2P9dtN82/KCgf646WzvJO4BDwnCZLQGIYnsOQyGaGIMHxGrKk4vA2ZnHxhLw180r3
of+DffyjML+n0kmTdYabKJLIOn7iOziz2Cbm49hi5H9fzBTc/9vKysK8QZBzGIfOckpT6V2w0fUA
KXq/QkDBlH3HDRvl1wXo9yoFRKL6us/eiNoZwhD+IAx0CxVAvbk856Kc7jUFsGdVRb1o6CHP3ehS
7fhkWHCYVXBedc8Yok2p0imvS/XF4xDEcieFTmlEmqH2QjO+MkqZiiBIS68TFty5f3mofmPFnx1N
2P0n6oS48MEEQB9uPetFJjE/jJus2fKQsUH0sVoNSeMR40f1MA9jgoEwU2o8PmMvrw3n1ZucNSvF
ow/co0JrzXB+3JKgTMUmn8s/4y90P12yfpiNHu+rBry1qKT7YIo7ye4o++thfVhsoLjjU73IznuP
lslhRC5nV4NNzRaChNEF882XJOcrRS2e3UPs6OSUQHuMFM0Mkp8ortHR5Vq/hB6QpYNllRdC4d/S
qKGk/r7IHYa2ibgTRTfa/M9OvHWeZS9Vw+iLe5XqwAxkNru86/XnGPoWloOV2jEogi7zYPF0+MAS
E27TQLhiuqhKlAKDY2CBxkJPYfTpxSJFZmVJZsw0+PZtnIs9mc6qGGxRRTFRnGfKS8IwMExuRRM5
b3jm1bF/xnevvADDmN62Zt/J6CRtpUpeC7Re/TtDQiP0l7Pi4+u83Prcxu+/cKChqdwbkFPALwKz
pDgLNNV8yNXlsWBSh2pzwaG9zxfLcgo/345Y397XSVJfFceZQP5u1X8a0M8JmcAxgg4sFGzmF4bd
zsjHK8L+2plLEocvdz+sRJHEPnjQuMtqWOtEEmXaON3ca2MJVkiQzwrJEwUF85RcNeGHRLs1Kmat
5cokb7Z924NT03F2Y4xkXY2/CfnneP8fDPyv6+esuTfdc4a8LFgEady2xI0ObXOx//HtRphJi/oc
H1P4guoi2uHe21wAbqphRlF5L/Bm+/QW5fkvOLjHyCY7H5ii0QVTuHhowG4pxz++QtxoKTLfLnzS
U4JQB9fvM7eAR9vSGTt0981JyQYm+muftJbPiKMbdEqZB8Gbe1sHlTXLP7ZjFatRuQgRladIWWPF
F/v6Sd3Ch4CVaQr2FFC3mG5NQRXV1CE7kydgHXdoBdzBrVu6QU/sf5TGlzf3jwuJVCDip8t5jo36
xGQEh+J6dxg7xjvM/HJlKCWRfEHc6Out+pVOPGoGXqRlS6uBlV/j3QvDK8x7HNqsO40UzLFV7VGB
+bJBrfetRkRv3jjPElYsSQyKIIFN1nHQVZYmm1UAmImZIQYW9ObqGKqCc6BqUhR/k8oA5DzwJKhl
VvVJ5fWrmuMkommBSkJyN/0aWyoIymDAYA9KFHc08E0EL25hVCINJ2SM2qM8ZSDZNB4vZ2Jgrt4V
D8VTXfsZCfSdTxUMlifX04AsHD8imgq+/Tq0xapasZz4uc7j00rUZfoRLJUyO5h+o8ov8mtPIK7R
EKKXXb9A/Dm8hr4/nzmZ7qW+sWe7LJPTD+Wjmu4JWPlIwf5Qs2JzSSLzE7E5WWhxBGIP+zcVgXwO
snE5I5rmxLYdzNwbI+S7jH5hXYlScRBjelPmZpo4e2K4rzuUzdr2JXt4APx1rB0zam/mRJ4eqSCp
a9yp3OhukdocAUaVzWr/dB7jd9t/0LfSbuZ5igc3tBwcSuDw3xbwiCi9Vlhp7/yf30N4IS69b4du
GZpuCYZMCoqjhqs2JVIWGVNeZTwhuysahYoeqgtoWY2pjbZvzgWzSJVoHru7OWr42MKDYpu95wlr
OKrL/kSnSAVAjIMqGnWo5iUHQ3zbNOlDqOMhDTmnfMCkL/Lmhq/lAmMtsfjuIfTSG8Xrm5FDCRG5
ssPMsQzcl8s8RpDDAe2GaQJmExWn1yGBB7na2Nr+Bc87+da+RnhJaVRKEFaikKAXsQksuX6yrNHJ
BpN1HYk5PrdTVxgVYR8d9c+eGmw2RrZFuayFplfuRWBzPp31+hxntVJwoMVhwxO0YY+ablEC0/Iz
vG8sgbgPdFRaJZI7JUDMkLVl6svMcyfLGrV+n0icBFzAkAi6husLaqgk/y6r9WlXzNL7d2IFUMFq
TMo+hsSYHYjJtEEy92hLOXAm9v8BkFepshaCwBOFd7HBWIG0Uo2E5M0BZT3CGV7kWTTY/71qtXYm
EJpNSFgMlECru+topNNjV+HexqCCu4JOAhJuuUyusRnWKZJTWdUNAq7RrlTA8IjDMxjv6OPSMwBq
w49wX4PQRZz24+Pe39jdysZXn8Yi+hCBO4e8jIOC2rpXnjvbBSDe/g3y8gop7VPlrGzzGYhV4y+1
W48rpK01xm591TM3H88skSbybe9o5Z9OYDGLiSlHPWghmr5nTMwmG+u0wE95NOF5T//7ziduaRrI
BJaBM86izuECvs2HppHtP7zS/qpfRv1j/5ISPaLK/p55vAvmp7WeL7tIwyTCQLTTbXFGCS+7lMip
D12n4rgnZqY0LiXzpVvO1v2VTFZHwYih2+/iVph2Pfcz5Z2MrcvGU/B3S19KN+pAPT0U46RxzHSX
Tz6DCkQeuqmBFaCzXlaAzdlCEJsj/ey4vRU3RgkpkH/1VxC9yi1LOQB7TOvs+2c5Q6qKbJGH1/f4
54WAV6wCUBydOxILEEb/wvZjzsbu7xbHFTV0hgSbXZXpsrGnUkup3WqCbVC+zvxJhXzoWGnTgCvK
O1MH1O31Bt7abd7uGX6JcMYE+P9JQCTSX+btNaAoD1uf6R/HUP44GAODxxnXoipXoF/S6veLkCJF
n9mJamBmfor3nF4lbKVllBk40vuWLTvS3Z6uZ9IORRAdUwVwOQSj9u1jtRjvU4xmf3VZk5UmJrR2
avz8Vgmciy+RPteif5Sm8D0tp+CQ1w9QtgCKhY1jV7lOiqjv1RuCmvPOVoUGLQpU3ouDAFRpXbTB
hfMY05jDhVJwivnkA6Pd4mwcGs4SK0uS1YozXtVBPqprcOkPKqe+U7MrMoi4liaPgCIcj9LPqKhS
La90dflgGIJK/6x/preD1H6KAVaruj60phM03iN3CLI/Qww8leJqu6bOS2N+cE1mJ0E+hSf+wHl/
vT+5POlFagNtX71/ZsuCNtoo82lnHltk2YJxkTDIe5fu8y5eYX7Hb5Z2V+IkfPL7xmpLL4d1pQvD
qoM2wDKy5G19mwIyizcTK7STXZOD8tbPHZZ4I3Hkzwgmdu5rkVuFjGFdyJvtTRhaD3JQ/0u0yX1p
YUwtcEOjPZQ/ljcOkoaeNYqBGYYtcrDXg2yv9wLtjOS2xOX66+KT/KCC95++UmTfE+VOTaAoh8AR
NGhLwYXBINs7XfkIHuNECm/TVXcvdFGNCo7eO+UdnIZkOcrcY2+1vQ+hsLfx0ushlPBA9GTdl4Lw
5AMFkyT+yoCyXFN5nugY78CDjorYnpKE/EMjTQKqHh3gRibbwzIcCqheD1nEReIENIZO2iI3aq/Z
Q0SPnDQ7gvxznMzjREoEcp8UnQPMckLrjxlvZ+VOp4SGuotJrcE/2OK/1VlpVYiWX0TP1uKcNa6b
DM9/RV0DGA/OrdY3XIyeVT+ZQdxKXl1b8UKpzKWWDq9Qtvr5pzGw4+H4zvT47xhRco8hDCmqnlR+
FuBjlfwfTQrI6QveMLWc9cpdlB3XpgZ32nYjGLxxsSg3sGLdIouEb/w67l9eXM6ObLWhlCct0SV9
gA954mZmMl1nERl735C0vG1zc0ecJEDsNekuiWriw8DoE7gRZs3yLczVantjd7QOqpnjo/FGNxcT
e67bGn6HpnW5Ioms8BC5+KwVoQcevOij9PqBYtFdcpfT94ad/97VrteSl/zaF/CqtIj1HX6sKyTW
ovTmFstbwk1r+ZumIQY8/s7gQTVGQptie/bCoUePqd2Sure4k7zIjC3v7ZzTQukp08adU1RrG3T+
iVyMa3zMOdHVQirLaoV4QdlkzUAri0L0YwrGhXOO4HwS+8muIfHIYNbmstKPfxsdqjziOzlZtP3z
QfoL2sPqzwA2dc5tq8aXRctHgmGB5MJydBvL1tFw2YjWQjU8pCI1p5i/nxv9vynt1vsDCSerCOBB
WzEgqMjAG5QV6RyMyAZpRAhpwMKFMBykOCCUcqo9J/VRX951bskd2nI62VCsU6cGaYCk+jSdLxzM
UVtXSwSgpNk5/lQcE79T+LwMeNXRKM95dNXUWlfRFFiSyqglBO/i8J4La4FgmiPKdDL+IQbGq95R
tdhdAbfHoQZoyjaeirsPe+Wedk+NiJ5mc9IAu688Q3BOavF+lLViNddD4gGl9xP5po7gBK+OLQwi
kte+nLZKVouH1Mfw3IgGgOpRSG8R6QalB8uW6To0WW+npO3A2rknAfVEV7bdcYs+bfN6Znoi2UyI
hNFxfIj9b5WrHYG2oiG+O45rAcXmAtO9noDDKmFmT/SgM4Ld01702qGZwhS8SQgaOiA+rh13erm4
VL8wBXzJbWCL7bhuVrHzpnVVNopwfmAhRpCgBwR/911JXyOZuwBO36kIoJ40Y0oAqtxGF2MUk34D
KX47AZUKGs9P7uMODb+pgZApysL/vZ7Xa4kVNoD0wVoJR0jQThgk4apo8QPUb2K7wafIdTL6ssp6
0SrcZCjlzkDkr4VJ8uzTyWpMtLVG+8+Hhu6jcp60r2c7FiIB0y1ec/f5b5dSgpIwfebER+tslpIg
vK8CAUJaT4prCi+JDASuAhez6kvtO9e7ALUXhRHRmO3aE9GmOHQmKo+rVmwJP6rZfxDbXahJQWXI
ApNA7FlTrIsUlvIAxrno82QfL4DQG4jhQCwUBg+Z2o+CVzTsdC/PHHbjLpqRQdPXxPYb7/9b1/UO
6A6zulG9belU+75tgRRIYrBB9mgIjf13hPxQPcPI27m47vuftkqpeVp8wXZKXqhnZkj6tqAVbwwz
oK1aN4uJWt83V3zzmpumHIEMZJ57XliE9pxpBPN7m2kp3buh8g6yWdHxCT0EoExXVQcm5YJ8nr6n
UuDVgEx+b+9HEmNxOVRFK4v3giPtdPUbusBaBiyhz+1OuVtnHkgUTGybyaZCUXYTYbCX8DXEBrXI
Wl1tTH8gh/WWJhd7iFNsS/fLJ+QjeHDc2vB7RWFDJVSPl4jp8S87nDdPPTtTpY2q3JPsOi5yQ4eB
5gt4NUbDdpLmYotBaXwtM9mpIayjtC8sXiCWlNF5lW5lW3UgreXat8PJQ9xUjrdBmOCuFsVIf/Z0
xlmMmwqbofpjb9ZK2pccywl0XQ48l+5m+HyMykagkggehUXvYE3wU/HWUbfmRK6quj6kvIB4c8YM
Hv9dOPSHC6u0zvLDarxGiVi66DsuZvvn7YTOcRbFGwSzq9411FWDHxh+s6qHNHkDALLyqIHuVNVd
ISH+Gr28RTK4MebqY3Hx7hjmF+mGJluam8t+0Ag5m4seA5JBq7eqTr3fg7I6b1TJuT3UkBgkpgxZ
ryMUUMRa4PcIx59m3wHTtF3zoovIBAUmkBYeLlPTujVRCI3dAKSu+cld4jamFwAfMHJH5nj/YYI8
t4qMikK0a8AG99AxZ4AmCc+vCVjXph7WnU09x1/wnk5ktaqx1znEJ+4141BjyP9t2F8Z8R1CNGZo
KJVyhNdw+I6mHDUGHAGN0X8D5wXaSLOs/ifzW7JFG2L0tr2O182WI7vnWWsnrWIgns3K2zTQMXSR
Xm8iD3Qzo0DJy1HI1QMnfJyugxO09WAk064Z9V8xAg67M2S6VeCtfCOg/dePTLaIh6jdm79nRnbg
buE0scQLicwhuflx8TeenVJxxOgOM7pdKG9lrTSV3hwFDoEg9GIAEckPlqdbCtgvflYNSE00WBHt
//hmfc2wya+/PSyS3RM25FxM9f6sgmczqYHNzdv9GBCJgVFyz064/0McT2GwHizt4IBxaM0cOtKs
dCAwo4LKq0jIotwRHsI7Wttb4Eu+0KS6objEbY0w/Y66crH9aHQrF/5TuukQpYaQIsS6wdDNr9tq
bQ525nCtZw5foX8Yzovil404UQXux8ZZdJAuoWj+D3dH7am1KIIm1A+OgGJhYe2LQe6T6Tlfto3E
NyrLgtjVBxqgch5Z5USBd+6KtlYyUcqKxaD5oFf6jZ9X+EInD2Syy+zXkszZ8lh2oBk70tpK4Mep
9OqOLzf+XrUC4W6YDLKhBeZvbTPSrnFaW/zBfZwlsXFgAWxGFmN+IkD3C3DxStibsrbwPO0/2kgd
ik9NOzcujBX+hzwJH/0ABnPRbaGpNfmTEoqujaLwk6aqqx8HlYThu3CxBvcmdLur5xdtDB+ClLca
07ue/N6gvSFrNW39xNox1BmNw4MskMaeQt67qymnJ4npyS5m06JTblcVd3P6lEse1E2aYJC/f2Wk
l4jUSyf0RK4OVkrpd1fQAxyYnxeaJCQEwrZjwsfnBoGSFHTjlqFZshWzav83px5F+GAxRYOWI36l
9ySXjtYxCj6WZqng00RnHDll4Uq1RFeeo8o1lQGvyV1i+tEaeRPW9EvK1zZQs0x/4DpxWv3LPfgU
OYq3RGaBcumaLjaFCxyOr3bxZzZ41svFQNDYPtHgiwp1/g1Q7p8AoOmZAvYJhGNqjcZQRuqo6ZuK
kjUzfOmJL6Y1eTtvkm2wkVXtYSa9gt82Q8zwb98TNY/tDGolYKlRxjqfpNK6qiDUO0sHk6xGlLrg
WNboSIpRXuRyjKiYD/Lmjh4aPkaljp2fvJXp8bMCY687QhF0WfF2rPzYntfnv49ouShK7MwHQBL/
AZQGFAduHeegaMZC/kzpdhUrSRTRBwQS+fKfvqO2FNaDxgn29TH5RuEae1mxdQ2hn4a9zTHowgnl
SLsu3Jh1IEP2lKdKe+GP4dM6q0xTipFt8llomAuI/yO1/tie2IKWt/etDQU0bOeRGdicrphkidNw
b/f1pIJd8FX9VOm6CAkbyLu3UIl94xBJuqqwbnye4uqRBFETXyrKKFPvGhCgavA+uLzYnwNG7d9i
A8MCQq6WXUh+Wofrd/Z1KoeRz3YALMbigfAVD1caigJRNFOcSdAOuiH0Lp3/0Ydc7M15zdwWMG1P
YiDimQBM1dfGhAB7EBvWRrxcIQVobXAvr6HdwxAyrDoVIXFAvvDk8FFZ0Qr7wCc2lN8p+N65V3KU
ulxr3aNOKXwPBCmnssKKJsz31zYq6cDQHRB0WLudIe+IjLFtT+hxsxf1v9nNNI5CxwmJAP8wOZsu
RhTsochfvRjk/A6Ignd5n6vmUmkAyKgQPPbV/Zdvr+YWyr0fFufzsJDJKdnc0D8ID049GMi6YIKq
xS9xZPxKc+UP4I+fszUCARRMDKcKv8gG1+X8/SYU9wV6STszsknHU8LbIC3gJBRVlnKLwxlFaPQh
XVCqKxMZbO0mu17ow5HrRrosDAplsyVbKgXFZQ4puUJnatrmmC7rZiY/yFH4l+wg7EfBZejMs1kx
spYRMILiooPySO8NLlxfIptmv8TzjZjWgDg2BlVczXyaKzMZP9Luc8A+iLxq11TVvBH2zQOTfC6S
BVWaERY0ID+bVE44ZwvxNvZWM9r+R78mZn13SlLOlbqcVwEPhGLhqmO3FFWH0xKUevaWSq8o6ORN
oVHTxg4sgXg+gShZ0ok1Fs3PWeUhf758lZRoFdI/gP3CiTFsvXwgi6xNjIFkLtC9WRHt80lmqfSv
7FPto2+1c42YdGggTiIdzAlNN1rRjiefGenU+TZ3JXSlMxbd798Pk8iK46juEGNTztJfvczSej81
QtTSwvzXnZ5x/y9r1LD4yz6+GflDheZROhOkeKf2D8QdDMgi9s6TU27E6A/Pn/DV7TM1rL/UCJ74
4wn+wQK/p8mrYxfNoYtRGYD2xLPJua104ddjbQx3swZUjfqEXDqq3BH5wljmjS11cNCUViCweVgM
TTd5hRkytVAyWKCZ4iC6yF5wuxm4gIblE0DZ/5iJLBjmkKAz1psqYoBF/AkTv2D+OjsEAVyHrcIP
7CyyTkSHdhQTzrBUB6gB7CVHXGVswmmpFoVf+9zWPQHL1nC+NpTJW4MuOpWQnj65UKNzdqa3Cxvg
kXlvDafQP2z3z38Cb5fRCCV1MP39c50hS1AZ9jurnFcdAMvrSThaLY744G3nFCFzXkEtdMSgIuen
YLah45lNkXIh9B4tNDbKqgMDhj3j5f927fZa8QzkVRFdJs57maQ3iLQk0so2Rql5TAS9V8UtJBVg
SAg6oBd418VJEPlyYTWs4ZJDmGPXKoDW5hOjdrqSDbDxvRqJCB9RlfdmLR7RACkeLIZN0q8kNiVV
qHdP5cCW8+hGbvfbOt8ocG8DjBj+ngfSBDkE1fvtx/TqSfYhITqw6lzOp8vX2vLJmgkyTLTMe2nL
Z14ViviQSCOdGHKJjp/RMOAWyM6d6DsVVuZhGT5CPzcfneskJAIsSJDgVGqVWFZv1/jSmcXzLjJv
g185vpOoJN0TSvU0KWWJ8QU2OYvH7VWhRQRG37OTsZmVSJfy12llsFTFW4UE70elquqiT/RijLc9
CoOTnExGUXqEbo+mVRTaAl61NNp+YJS6JDkBeUhLfZHM8dTa7oTR4wTYCeN/hpSWmK9gMUsbvBpX
+RdbH7s32jYFlowUoUkr1skZrmMaRrePzqcQD9du6X06M7OHRDhPdL6V1Ix7QPrp/TfDyLsT56Bz
+9T7sLXHohwKt1CdQXubJxCPSUZLEXElCHO8Ypbuz/Fy7NYXruedztveqvb4ZZEC6GTR8gEkfPNR
WyzlUII2zsEdp0mLQ6TV5I4FLjehbxlw6OBS+a/BcTfmnm9rYiYWBUXVr6a37cq8RoUF2atgaMvV
5r/J6Wxv0NAC6exCkdjOV7XiyM1lIV8NTMbD9SgzZLvUiTuVmaV+ZyCVNBCDWVyRFZzjfigs5TQY
OkRYL46OmpoTjZEe8YcktOlEX+Mcht9IsOkr/KreMi7vib7RbHMfR7Qo2AnmRRrMe49gHie74TuY
HHLqcIWLwrlkfDurhndmVH/UWRdNLSesJizlV4Qn1xyY2Z+24pghMJ8E8WX9GtmRDcH/1Hi+p2ZO
r07OMwKi5jmxL5rkcJZt/99C0iyIDhHCtk+FTH0lrgFrmwwr8N4mlnnjwloyJT3NnUtb8aYrtk6F
aKtjivkGDP2iAjVvARjEJ4ph23/6SNSwtf/YXRKZYF4q1cq4ks6IsWHuvV+PuAQqyCwjdeFU/rqP
E3bQLYARnxezFixLllYhLL0LWfD9gPRlYhTrKg6i+16EDKTTUfl83mfgisSvrjOqsiB9ZSjTWKLB
n1ozp52pAY77rFkW/leZrobVYVMG/SpEBmWDIwdWqo8vSv0XOOQc1O905LuZtIMJDlyyoh8ab0VN
xwkVY/akd5AYB7v8WJ6fB+SosXleKPLDEdo1z9AK90IPfUTdxCmaTlEBUi65i+Qcz6+MKDGsEJU1
KkB6ytTLP3iIP6z/73gvTLBH0ygBLSZHp8CCvsyhJHAUszxsz/d7bczt4o1mbiHpkvJJjiAudt2K
Oi9OOm4vI3x6DyL/1KwwOKX7RylM8fJqQ7bRX+sXo1819pGiZ2gK2RcLQr/60b0fbYCBp36MKDAm
chbYUvenNzKRDljzOE3qhAJK/+H9InxiAsDstJpqyVrd8FAB1pd2UsnCRNnYB9LB9/PorVGt44vV
3ZD57RlGy83AGTtUyJF8J/x/7Tyb9t5T7QVoQpQIjc/U/pMgBxRcVi4qvJKF85k82HfnjjSVMquO
7qEYWn2FJPcF/NXMHzX4sHrQR6AG7wq9/nzmq+xJRrQ02oJDTBMK43VfFRnfrICIF5gsF8mD5EJ9
1otySBe1IZN9w/M+F1G7MqDHDcBnCJVc/wbRCJKyJr7PuEdJj68/OKQrtqmlMT35c6S5Czt5ITSE
zqGybiHtd6VXnBRULxUE4meWwgfc64GYN6EVC10+dGIeh3d9s81s0OFv0fP6LXuNBlvxFBmPRSCi
BSCuMtk7oo7xtDQd54FL4Vix9pQ6yjts1SULB4CS/vvWF7n71GF7/8h4U28xnC8/YHWYSPrBtxtZ
JpOhGRZTpzJfahvZF7UYyLQi9XuvBxN9yjI2O/uabcrUqDtNvPjrr4Hj4m/fx/XE4HU+wSpzQL9E
pKVzqcUSTwfr/7K54HogWAmpgaDze9LRs4qgsYcGUYUktNEqBQcOZDWKAjANkFMRBOjXJ5/t/MRV
UQUiJowsIM3Gvcn1ySa5dXqKI08xe8RddVxy7p0Dg9nqTK6s6w8RgSQLHJMkHl3ZY5AfYnaJQJF2
OoXt5gZjcRELOVSteRz2weBr22kfEex0qdVXxwK/G55x1dUpz/s5ll90OnKtVeFEz/c8Etf+9Wbi
k/WKDy2kHUlESbopqHkVJKish1By5fRA68QwN9y6/bqUo3JqgkiZvq9H0+QyUWOAw5vPA9jGBjbE
85sGs7KeKENvz93Q+lbQ0Z/gBq1O+WpYio7oWb7yv4ZnTzc35tawukAS3xEnzZTMGmqIox0VIGxv
GllEGaBUfTkS/IzOid9htqxmbORnS9+e8l/THdzLBmRbWxNMje2uY8WNQfXezD1bR7cYPEiXPw+L
0Uk2LaigKbiNbyDpJUS+kjXHfzj4XxjUf2I/k7vr124o3ktOufZaqwAiTr0YlVsdxwF67q4MElUH
fpAKFqxURxYgYiWsZ+KgXxwjGM4uLZeofq7HDUkB81jeCEyfuCq0BnqbHP2nTOpNLhKsCJ3lutbE
oxwndMHngc8It2XVfmLNBVnDJlTUYJJTq/1vxpgdRAzXqlYnY7u0/sYrtTMq0wx15tDOPS17/R8y
a9LqhN24QsC9C/0noMk+7Q/x3yIbm81ixGqcH8WS7kYA5nm6A01DYkgI1lYZP0c9beZA3eCXAxyT
+oct7xHsVtZeHqPM8Sv8g0dATUaNkpxq4cY/zCBaSCs+I7oxzz/4I/mk60Edf5PRTF2oku2Gwhh2
WSbckzCvMQVP8myQbpDhZOyqRTduPptFbtpjla1PPNX2Y47kq42k3CCy/OW63yDZ41Itif4gGBcP
iKCDP1y1imXFeo6s8mDkM4fnDt3yb7sl0Xa6qlhmdZ7oEdAnWb4HebpuuT2LKdooPMVn+Bs+sO/d
91tNxkdNM3drLRBCqK0e/fXg/sChJ2B5ysSxEebeQ2bxQ+uE7I0sRSu2uMROPjN3j2VSt8D0Pdhj
iD9EtxL3XJtHhs70lh7xWzKmuKqkTmhkCmxwF5SOR6FWuRmQleHj2admSSMpqg0VmiX91MwyKuEb
bX1dhC7YnwAgFom9av5yMK0Sc4VXLDEgipyQ9ZpCm60ccOmgDYsACayQCKTDIlDqAK273oe7NWyU
8q5jlCB3sCI+ZzT6ovTN1B8CbTX0N0OigXptY+7l3imCfGNHnrEWuvgCa6X4UbjlAcozsZWOMAi/
SDFC8vocX35fahfjdN2O/Wx8pFBjmyzU7h5J3h/gtd7S+GxDwen0sP+4oM3alXYGXuliUAT8ePaB
x8IjWKr3ispP49/eMifpgcY/gysy4ZjDfYgBY0CKHgmPjwrnDSTw7//udjkR2HN1ZXKpbOLfmDtb
sEvQF0y24y91rQLgrH0pEpF7Q/rsTYc95xLdaMzSEkzh8V9qyqubuSSEx8B9uusdaE6rLWzj29RE
yzAXUuFgxvKm4zX9tgaVATNGkkfXv/D0xTYsicXzRt0inBYWMf5gcBfdXpspXgg5hEzRMOp/wbqC
3fEJVeKOtkNhcIZxlpTFCCwyVl237LvTUbT5Az3+DMGhNy0kGn1TfInlJJ/Y+Vc4dhJdY3Q9wgvB
r4lhj9Grth71zlgT8riR+1U1hXKpIkiJdOTILUrH+oi1P03i/kdvcvg2GbMk2YOrEsM7YtkfYhLd
4g6SLZm2OMq9oucYnMGuHy4+Aesunfey9a6G9BLefq3NZ8K3viU83/oGfQrynX40Q503Zah1ChJX
zWD4jjSeFMZZsywf+exwr3zHEw8F5dZ7Zn07qklhqrd5xrXTy50dzDzQlRkT8jyVSODXGZ/XoDV8
FyIR4l8R3vbQCByaDE7TbkdKjLGQoP/BTEoqU8bL8R3uhuzxysOCs+o95EtSJ2ONAaKBkIt7ipEo
0FghWMQfQIwbM58ayOSVITTFb2bZeSaySFTcLPKDQWIWelumzJI6V2QRffujMK6K4scZu4g1JT1F
SyEZOR0Nc0yaLpHnoMUSpTObkNxBNmbxfzPdtIaOE3GVSM8w7sb/ja1ItiU6bQAT+xqM2j90iPyY
k5ty2KOM5jra36YoY++85ioveUEXaHcw2iMYNqcjVN1g4mefGzIwbE1gFo6tzprUYnGQB/Inye3g
szomMZqoDQlPiAih6iqcMKrsJ5MT270XGqyL2Cmt8XUf8SoXhzA638S/3OiUvpLk7n0aVZZmVj/v
m0zSvdlqu3561qW0DqArjqH8UDVghKTOTtD51h1VonnUq6WhGQC9JlCbQTHlw6AEJIIZWQx5YbLR
zH2NKWsL+fYSB4iuLxEom82ivIXG9C4U9I4TBZQ8bAZyLcV3CudmfWgy7elRG8uLG1lqA+LOWQgt
3SwxEWeAajYhF+Z/MmmnlOBVdsYalTaQMxtKZfolp9HbUWGeeX8IM4d6MElajGHIdAlFoFMjcbcO
BVbJOw/y/5xMfMe0iG+Tr5k+oIX3b+Ul4qo1z+znJy9l2k6tj1v0yRaO6VagisGZuxvpl5q/4bwL
QbDUP5lhGT6LkGWCfdmn40p8g4it3OcYp3bBC7QhFQcL6NIqLAlg++A5vX2ifNMCLb/3+2JQiSIv
x6uYaTRXYt8Jr6tiZX6xKqd79P0uRqAWy70akUyyQmQAFTXXI3HV4yDz2P/UTylfJlOy4ARSFmd6
8XOpWncy77REuBncF/KrBqRO5M47qkpKOWm5AZKfdZrSCC84uVrYITyqnRiGApeQR3/mXTlg8jjx
Uy62tuETq2ilFObQ6f3RZJFmjh39dANAf4+kDCqUbxcEzqHxDkh0j23wEfgg+r8tZhTQmRz5yTKu
U1+szfaeqgxzHaXvgKcXm+esiCUDLRlpfvBXuSUMyfU6mL3AhknsrNdCftbfaFR+shDarEKLvrPw
H551NnG/WCeSqrTRHdCdBrH1db+jgKwZvPqHfZHiuKntotD5EfX55UmkzjNcgMPw9gtdIKuNySPO
Z33+ibe6MxSWVBE8QyW1BFS4mFDCMVWN7Q71z+H77J/YjGQTHVzmdHs+Iw/s5m7D8fvFEMtxY09n
VVNsy9jzIsFE71FXWzwqAHpPkcOyDV902/va5PhvaBAKK2MZHqgXnpsVNlmUi/c/+8XoAS7uNA6F
xw3XaxmjIw4n5YQcv89W0XDLY48xpHWJBp0SnOG6/x5qV5tJpbG2VnIn14inTR0GnpRuGhJnBuDt
5zr3SjZ7O0p4jSmwpIz8ClvCNeFEnv8xqaufCBrG9uI5kuAW0BtAEE40FXGzIkE3iLjWheTL/LBL
tK8AX6VrSJAOfNNu3mheMZjNJxk2KkWhMUlph7fyDFxi/7CoLhG5dnZ5NvYKuKIoU0xk5SD48O6h
EjivyKL2XIoGonf5+8UEz77LjGdl3b0VrBlCowBAI7If0efKNrfKZaa6znjaj+8zwAByBMVDTnsS
/sv1cpDVe/ZvhioAQALC72UB3lLySfF01WXjk/vDHsZDX2iMhKB6kxiflg6roilINdU1yvjISNn4
Y0JrZAF0WgMA7QWLkGn+v72tYCyhIILoyRMkXJJqMPdLRtjLy3bjyU4Yo86570kPiNd0WZsBo/wa
CR4TzKkDl6d4E1S5hx8oZApmpSbu+1HtfPp+v8GimaI2lh+qEHwGsWvE9AivmflDlI7AjVTQCd6O
xS3lz9KkUK00XBexU538vyJ7UU406+w4uVBp/yI1H8E19y1HFmOZTcvO4gANU9/e3lEzQripp6zO
+xQDPALU22BIHKKwO4hQtP9PonbWZZ4KZxIHsPlkjQE67xg9WuGIThSHA5wK+YkWayM6OwHbPuOU
ykq3Pl3HCPMY+coChkYTAxUGs/kZFbt2+p3PC6UENhXBMIqZZq/wLT3ydHVBkWtaxrmKmk94OcnM
NkD58Yg+Z8l3vAIrttWTjH72gsMCteOZN7INuenBCC4T382lWUDTmvUxHruwcMhAATNK6b6XYorS
8W/Mbk1zYjT8wTICiPVY1UlxDpzeFfpp10YKv361fXGtFZ5ahpOEsFi6TEucqT/xHOxfrxZgBvuk
U00ags531bqduNGWgIKza5EkzbQgbTPuMIRNeiM8feh9yX/nRaYL21jywPM4WfDQBZlW+0xuHeqL
RvW2ASFl1ELJz54qWajCjgA+EV9i+2tYuclGAWULYQbcK88Lei7aS2fEIDfgInC0wEOI5ipxK7m2
vSE7beoMmukREw4Dqs4inFJ3iXC9wxb3XqS5WPPYgSWqOo7BxH92lpZKoRt3veGgtkxVXrEhfp4H
fdaRJ3nPys7lICNFneZ6cVVoBcaHh3Cn7k1KjFtOcJ9paW3UTXNvfDmoM8ALcaI5Sn/ok5zT/Jcg
Yi3Jqp63RX3MZkrWJ5nFEUrUaOCycTUs8cJqAtHjnhTJrwZ8ned/mHY7DayWTdTX/7F4qLt2/I5m
acV6xxslZtaez9keR8aAkkTrDmGrt46u4L10QuxRAjeCjILnBjeFNDj7INKleJcHrIxhgtD6n8EA
Jk6q3MFNKWqjCxqE+SJSUVkb4eut9bMqQBV0Z/y+4N80O8RuKvSbyAkecF89W1qp9Y2iiD6iRqbn
BJbaEwjiHx/5+wJCqL2TYsr9J/5IEvOLoFRKSt0koa0zK1OPOJkwifBQyJ1vGjsiBsq2fE51PPu0
VySIWAI+d838u8exEacvvmMAysUkwQVFlq5gtnmGvd0viydiIVNuiUqbx7xcmxKotpZkdMgLd1s8
i+Wy2VmrYvMe+Z2Zf6kSNjMUkzc2jK10BDd/T+McpW4OYGRmd0veLyR6aWr2PVuTuWr3HSL82kcA
FMvIe3YOwx0H74Tm2v224eFwk8D2uUdYXPFcEl6wktmWDuOyq6ZJyb25llAdP7qtKgYxGrG/YEnk
nMhQbYfG03QaRhIwkUbuC/dtqbpUmkJ9H069jSctkTrku2co+hy1xzn7wTqLXpFtvx3pRagRkiD0
zPJRphLAe4jo3jchP9FTSeo5sCzgLbpBKN0HZnKQVPFmEEN3fPY0V29afXIjmVIzR9UQqrPT/ooh
MfAt+EO68B+QGy+aeoig+GMef4eEbvVBb6x9cLMkUnPEs2kywjL9eeTId+DzKPqQ+crHGSU46DX6
GX7JsTG+YK4JFZWFq1yuRdP/P9nLWShp+3YSaFHmNL+oXR4DPdx47wuEjsPIfIIMzoStIAgwURPl
NNVj4HUhxm7G3AjXAkAzSjhPCQFPYxmYGfZTU+MX2dwN9CZ2VefG5OI1aiNChYG+JtgBc+pb5Au/
pD6WDbLPCI8MyO0Oq/RE1XedM5PhcwtteqDfAou4bPolwyNBwNIc8lktARDjeQZGqC47Kt43jPYV
m6coLCtBiq/CC4SXbGS9fe1AG1nSqdWg8TGgGcVTdyUoPSPL332/obU/tRDMAyyopA3WP69HpVHr
Ma+HiT6MoROQeKcDwbC7WidN8UmwwasUIgKOF77JZd5dIofL9Ou/yOyI7aaDeBrLmrOSu9yx/E5t
xUnd58G3emsLXexCsrtqVPOX68a1N4JEEvcg22ke0vkoklj7epx2wn5VGh6qVZicpPu9Bl3Hojin
4g+3/KRMspfZh604m13d3MKVwMJ1qe1s+KJxhqge9LKBZx/xTXndmpt4JXZCeCgKExO/U0977Gko
1qvoYKDIh7+2zyPjh2/9qnUxBC2IFX0EsHfCIx3bKQvKpJiSr/utQB3pkNEe1tKtyskmvsTlOXsp
tMgU30ut2XMoSp0ecx9dfed78IIbuheu2PwW9sD+Xmd5H2oXVp7SYZpYMRHipAa2dC/PZ8hN9RR/
NdwEV2G/JA3DnVeaPrS8LAUZcOUl6CaSea9R6kw93d+n+uE4dyzKB6uYeWCgPFnqVWVPbJmwLTHY
MT6MLedr2nC9bSGBZ40D6DbCeZHa75l/3ZJj/26Ued43ki6GMmhRBzoZbTMvKipS1gGjQIv6yXE5
z2h5UXrL7YqCcqKY8RIESn1sqIY6ud08/5ASfz96MgeXI/ost215pN7SjwJceh7IExQms6f5rvAV
ZMq9nIPIHWcGCRFRf7QwPv+VHxRosTYLnAEOjmhB5ZDlVxUJBgeZ38Jd1MqjsfHMamrRAzibctMQ
+tGpud9F3QiCDARaCE5IWBh1XaMoLgH5hpFn7m0saJIYZpWDjQkjePtC+GEux4QnPsZ9eRfPW9w1
pIarFnwGVDyfwLMubbZ58mb2zS9X9Xj6SZSG5ExtZVKnmbhmxTsZ3wZ6YCZAAmDBUJSDsx/eu1in
LZ6zd87uzURvAVP6DbqwPyvDRFVK1qx/1wYsisLtKplX9ZJ58avK9rwYncIDgZS2w5O+W2rf8zEn
IIAHmpEZL4sLcUwXLUiElr4Z6Iet3/tHu7Cx1z+Z3tsqEbBrYvyN8R9EqKhCxNlRWUAtXh8EhdLx
Y1gf1SRjTg/dIVEkwEue4Cnsgd8oOTAjxa8Rr0YjEj04/wgVXnX2EFRdCx6ogAXtdiEaiWc5pU3C
EgyjlJsudFbZ1oH7WyCgli+qQI6mqZNgXsSai0hwxOSxnL7DD5VKwax73CP/k0IUMsYCsf4jneBz
d/KLRpEgdYqu6nmdveMtIfCKQeZFycKRo/IANFwZcUxxu6pBAZ4iPh1RgZnBNyV2CLPQkI6c/anT
UV9y3qbzf3lCVY+62zXwgL2PlgozRku2Qq4nslX0cYvADPAELwa/2keKyUUFyzWVpdPV/zcYB7qN
sRUE/l50e2mDTGvXgTNgLs91X2o6ACPLUVkOb9w8htzgQ+GIJuv4yE1NMfQUPDAnBMhdruZ17P42
VedC02WxZJYVw6vTJO/hOUCFNJIzcxWHVk6aNYmpDRMa5e5ICfb8osocJM2DVoUkU9CrB7IjVWz4
CPNbE32FsdScOUwqQlSANjQGZuzg/gxaVjj+B/jyDUaJ1TJOon5eamnxsQfifVnNXj5KcnqR8vZY
KP3VhJe2WhNQtoQatLovYFQT9n9KhZ/ZYQuzK6IeY2o2CvwEtQsPthAkd5hMYKtT+z/zEISwxDUC
Tx0f6oXq2Jd/or0gNsN6l9DHLmfX1Sn7IklwSoyYobhj1Bc3wzgxhddz55/wEGuSvvLM/ODMjJO5
kU1AGeU0cxscE+cYfc02F3KY/p+cDJBOZmoUdNcUKhnvazkI0WcxMGAjlxo3kJlPgxWC1iJQL2AM
5nTZUK+yFDPG9q8QVqomfCtjXy9ptL309ZUMn9X7bgtX41WwFcP3PmmKYk7YScKXhyxfWrxw/MYP
DSlK6sx1FpWEA2hxa+qQj35IVwGzDckuFCGLe3ZvgkiGChtW905LWl6BXG4uB6VEs4AI00g065dX
qHZBB5c8l/GDNA6H3Z8wr5K8maswOVCvY1wmA/Vh8vyjpCiDtSzYXTLLcNp44gOBRDDTNLvCPi7j
OHrqqtFDNfwkDM6bRbNgodlw8hsHKXDhor7uEjH8wX/tJ60CvNeVakoOcAhC1lTLUUEatR42uK37
w4OTpFw7xnbZNI17WF0hxZl7QVOa2uN1zhfEmwV7MfNpupNlDwd27rAwgxjlX4kMuRSnwDCTOe/y
b/LzkGlBFRnfWw7WwCd6cReRWh/fQzE884078FO/X73oihHDn4OeYCx3kODKY6aRDqRZiXCUYIIs
tRRo0pk0L+rR7Yy7oCafcqWMgoxuaZyDtqS1xWNpeEUr31mRziPzDfERgWbgn2PrxirxC2a/7uRl
NZkmgE1wTioh2O93cIDYu+6nOo7YSeh/dsdtFLek/xZ8D36cR5tJfXzMHllew9yAz9AxeQpk8enI
zUHD+vviKWRT4M2xfRSBvGnNxDrPXGh01yFkKg0TqT1UW/FTJ6W1JgClTLOcmtwf2sQHou8D8sr7
QLe8yigcqTBc6PrJDjYXdbRYLDFLjLUkZvDU3FK+9ThkCtR0rpm22m9xRysjry3yi0qn7Tg2uscG
ATip+cjB6FvD2mQHOdbztvK6cfxskt+KZJMexiyo6utRQiPtblaaDSqt68/aVL8I2O+AdwTDfQzf
xT+TiCN5dmX/sFP4nXCMiv9OO0WoPvJZbrNwhBhPyjQVJv0eHA5F7A/UhKNed/0W9dlLv192IMgo
hntyQ9mfmIL2+XxRkglRaCAIedxSKNlVxcm6MqjXLqeAoWt5992tQSBr8i/3f+KC2CWkYmkEF2mA
4wM1SC9KoVAN+NyZwI/s0Smj6kL0YiFF5pM/ZXDHSsOwgg+aCOL0LW678s3SzO3NSkzlrSDjc3Wl
RV6Uk2w7kku7NwIps/f5K5ijvayvZJpmp9Kjq/kgC18SF3kU+7lFiVdghKgH/ccDE/nuP73c9uoM
4crPvQ9Rleav9p77o6e6vLlanjBkNlImb1Gl8y4kXlNkrLYxMQbJZ5yhlvjmgM7WScU/4Gt73/jW
ejiRX1owKwtzqJx5g9i5537xuha42DrujMQuTUy5pT0tr0vlS15zlqd6vasITIaHv6ZIsNB2UbyF
AH6jbps+m4T4fgTUGp0eVoP9VXsbRMc5e0MI1jhtGrZTgtC8gnm6lG876/GpyPmh+0IHnwVspjhi
RBPyh6AF8ZY/HQTmmVDkv8luFM9zRQO5cpKdjl9ZupHnjqjrA4tB6t2COUac0EcAsOd3Y1BCo1gV
+l1z9nTArKfoUoNtG+XSgAHBf5hdK2vFgyk52caqQfw9NgVVGcBjbMdsOVZr64h6iUoTpdXEojY6
TACV+C2KASVLhMWf/T9YEE3P3A/U73f1aR5BafhEIxVCZhK5FXezfISDvYXr5zgkEIl/x+dZKSix
JLj86pHOIV7zKK0T326UAU7b95da62rlTdX8N/l+3YC9IUdeulPeQlFoHy+z2EsXsVvPPJZYheoP
Z/2PJXWxcfWc8G/Ve9muu5eQMNIdBCBYs5Rhcx1SOI3Y1sQ6bOzR4Lj8vXwa0duwKk313XKx1TLk
at5QeWmkHm3OYVbz3v0oyBx4HIsywZadFGOZXvn4TGfRhxXkOH4ku4flJw7G/djotqJeu+jBvhZ0
B1Ero5TCpnba56VblxAXTw+8o7oFH54cTAHMfWPZiL/OfAeFPdc8Ez5k20VGv8SORosOO9tWCu/7
kq8tyeZ/zFNhlsSMw664wLieyFGDHz3cShXmGbDsbfMoWE3jHHraQDHG8yE010f1cxn+j5sCaayY
HvIGkkh4d5yQhSaNJRg3gjilT/3cOQfQ9mtwtTafs9cu5lfZczWdA8stOyyBOM6QYcmM1RmDfJCu
wJt6Zk3yCtJiNznw3JdFO/e0hgMFcRaXbEFh6OBG7T4MtzrF+AjYEK2Xqr9UF2sDbK2nVYhFUS+W
C6b9bS4r9aII9/Wfg4p7HE8Ih1rS6jLIDwR0s8pYPphJ4G2mwSWTpkqSkXQYUbf6t+MeGWF3BCsa
n7oLPmAbq16wg+iVkTaiOFA7/vCTvEpjKcdaZT717TuKMWxoKaXcFYeK8Ko4hI7BLBiEATWISpxL
d1JPPoDXcb9fOUJ4QRU3RO/SvVuPhaC6yL9bbrlVB8OCuAN/id+WZ+74aoECWIqXyuNqS0WwzuZG
JtiZvZBueK8K+E8QiHzQgzIiPhK1xu/RXM6lcPPlHylnSxpFYgZio2AH6cWyG61W5h4Z+0JlCjQK
2bJEd+qXmOUUOTn3ACLW7F5He0VPH/uO23sEcLYWpGXQ3Fj/MTdBQ3bp9paxdEHCtd0H7niceP/s
ucYbKdDYIh2fzwLYCNP99jq6AGwHXAXatRhh3aal83lYHPHtG2LYI/miefu9xL/q41rDzhaJstDf
AgWTYcQhd2ZI4a6QLIKMbXkekELynlMuaCNbwaAapI3ZtyrrIjOYQQjZtg7Uaeyczqznh87MZLxS
IG2Hcb6b9n3pI5xaJ8/KdVaudUPHDCvAjyFKFr6RkvPvIdlofiZbg5nMo5Ksv4m6ikQRCz+pYcQe
KVaucDUUwgLNrmagkUcsvnL/zjEBW8NUNb9RVZZbRLGhifKI+O2LY2Q7t89r0CmC9bCuFAEfPxNp
pRhjAKCkCFcpy3/Urrmqd90mMxZEJb5y1c5oI/9Ci9UFCqaXV/d4pg0HmnYwOz0tkWI3boaBY+3P
RUV23zpgFxPBx5+x1u91gbcZ28/ev3+s14F/S89Tnt3ARS7su5AN8WTqBSuY3H+o4yu1VzFKjVlL
DtXESm50QgeAwiVbZPwQmLEaMFYOMotVhzUdbHRPPXySJT01YFeo+mFauKy39NIxiPZ5WA36Tl8U
IhWK6Ri+C5U6YsuO8gyVOJV61p/JsMsOUCPWNZtmxMcOn0ZkuyL7czErTPDBNEKWXu7K60d1JEfN
gDCONJVNkAEZEqzB8M1yoGcBvQ0VWeYBKTyfCwuZDirKljvO8NyyCoeef48Jr7lcrqNxxJmojB1S
EsM3ZWAeFbgST6e/sZiI5dnvKa7gS/g7P7VB/IPzpmc00AChsZOghJDp3sE2ywhcRQp7dhzayr7I
KyCXiF/121cmVBKTUVcnSAivrPFfOLvoNtGK8usPRsGX5SOiYBwlSMZaEZFWj1ZDdQN9/gunXDS3
ke/ifDeQ3C1okzOlrzFUff2IFiDr5LGRfT+PuJh4bXsYMvnJoDkyBU4qZGP0FCvL0d5q2dCe9fGR
LZLkJ5CZ05y1gqJh9zuJGotaMCfEWxizgFvDoT2i8FYQxNymClAs7F15GR+A21KcCKws0kdUTY8f
ALhRM6RDd6alDIkTBL5P4MdOF97mAK4mOXc3/76PeA9Gy6M+0TlYCrTzo21pS+nO6zK92MbQv5d9
ix5BTSPjuh10j7rtkcnoKZDpSxNSeeDB1NhEln6DGoBptSSz9Qav79pULpqZ5LtqTUNLyS3+jBk0
/czFZWf1Yj1ofNrS2SOkKslyZBkUaSIfxL7X/oNO6AU6a16KZUHPYbXNRe6FI4ilfWno4Hl9B4aU
Xvz4cC+do3igkYS2042lz9HiD5LaPh3UxuPbnDe/Z6CyaEokp5ACYhXgrmD4Vg9ZZQyfzHcdgKCp
dOUn7aQUKkJLYB55mgqjegb9puesdIpKYvRl+GyeQflnmu3432I+ZgBX8Mdp8Qz8rNRFrNmNhpAH
73MpdiZUlf+W9WmP26qkRTtIa7Inwun5+mXUMmsoJsVmAqGFpNF0gHXxUSXAcueXiL/9DOEwNAtL
5YxkWIL8ex6zFCQHGme8h2No1S5H1tzow2VlG7/LADOAN3T49Ffvqv4Bcni9Vebyj4DEmUQwPMaF
Z43J3/wqQyTSx16SyAOsreUVeCYyJzFTxD3diYnaKIX/9zbkq0H//x9/rg/TrBlYsW0mXBdkJTKc
DYgQOojXu72DvoYCfgocTwSnZ5botkTcmiGqynqE8drPrQVvi9tmtX1zcUalTxd1IvTRBJnW9wDl
mW2nlCLk5XZzciVsU1pNn9+GcHvmZ8IlHt8HGI753kcQJEDpHEliMmDVCo/YRZ36oThSELzbDnD/
E2UFhWu9y5DUWLPuwd7+bI6RnOUctaw7aPtQA7tfH+zxeJoGYOA5UUW6jbxeMmYkvgRWxFh8V/vW
r2MplpEOeKuJrLd0dl5uGlOnFwnJNTVuF8jqdVmAZmCrPZLlIsNeWCyUigklsBAkMkmuqobOE5fQ
SD9IACiqqXTAReeEkhD/2OVnpTVigee9PT5Vs8LOH/fUVZWaz/TArboMljXR52sJZe++KSFyxMc3
nnT4/S7T2L2yBJIxlzgaotfQjBtmkxApH900pFjT+fpg76lUVGyZ9h9Fkq9whlgCW7DjqXXmvtdj
hAgwU46wv1WUk9Y6nO/6mANzQPuZyr5z26HnFWGS9dWMNEoP9zFNQSq+c0cBfgyAkMncExTNROri
jb24//yjstfK5kCOGxyqJgUBnuDH5boo/cbq5Bd7+O1PDf2nUC23VPdaFILMvB0XH5abMiF129Ct
VnbBCQ37uEN4v6pUIccCQ/9uFI+kZ7Emcnm2HreLVALubEKb3EIg5TVHr39RuOjQy96FSCTuMIIE
Zvs5vMTABXnM23y2D2JfnUfFLSrDqHdy8nMKDVf8QbgcfyQkJ+OB1abPawwUsUHfrTHiIkuHYo2v
hBKC9RRN4wt+cLtKCnUPOIfCBCEwO51PFxWH83g7wMuUfWjrlgTW/Vk55GyAr0RJtzmNR79D1N4k
5c4Qo07+s/z3RUuHHJ2+LLkdA139/Ty8vcZFn+hWo8zI/RSIqWKlPxfVqZRahf3GzhRWKmYYBJe8
Alv5n5z6VovSm1Vyh9nuenPX7KIXkU6bqx0Wrxp+pFxzpuHh8PdwVRkn0uwpNmmcQJL3JKOAxIF0
jrDoQ4ef10oxH78Qof2PfzQGP4XBeh4OJUZUbvqRLbwLqTZO9bdIU1s8BeWPH3HFTkvBDcDsM3Ab
n6SZlTAwgVDOMP8uit6b25R73fok9F5hLw3vrFho2ZFH1N0jAnwhPepnNtPqIXMDinDCcSojgLEP
AbpmjRyePEPt9G0XXpgHxqlqobIOAUqFt1RDhYpagUwn4tpLa0fGfnEKS4ePJoNxzChzkn6QdAeI
aqvxpQ3hT4TLrEFZ1bZuNkahTWQWulQfEgBZ9YSWzKVQxFlswRRoobwnCKjKEhtOJtf6WRVombLh
twVUelfGo9TXLJmugdaLLDhUkpxjgxxRvEKHMPZwOyUm1xMpzFQnO2oRPilLqyegB4zPVKfoCFb2
BdYeCsZvKI+3AKIloDP1x88/O4mW/CkaqW7IVlxp6X7JrGxACaEs5SIzJ1FikGx2HXJCd3wxxgx8
uzSYf8oeYFOGZUY7podmmrUZxHOzQRwrSGyxfdcCBxCmJvwS6J/ylnzydVNr2eGRiGra1HGqekyr
94MXtM8QjYpjfXGlzI/X70Hx3KphYFLaM30fILtOihtcqP0B+1+LVb8hrXj2Oeg9+ZdgZT74Lj6k
9AnL8OWy42sPWpb5XflghhSTP89yMzeqZsnYiaibQOo5zpOsZmEmcjgVO2TmlgDgvwvlDsl09F+Z
h5Mnv2+VscrUWelagyNONaRVySnzsdA462K+cZ1G/P3UJeLE31/wpsKhxE5FojWvoI8H2lF6Gx1N
YELjA3UaE5rM86jDpDLgvqipVFZm9lN1Ul+VI/22te9avwpRnUWp2s+4Gw9+cxp+Mxa5EvXZbYT6
VCHDfzf588Ckc40IM3PDHkgImHzJbYA1nDzcjZe7QxW/0wtHmX06fD8KZ3VSt77QhTGK3yRtj3/F
rxEoB4dvyLwiZzum06WaCTx8scf1xEtSKkpY/1fixkw0vjWOCQEAhpgaa3vYbnngKsde53iVnlaC
QvK94siOhQsU4dXh1m0XurInqI0B50LEsLEKwZHBYLiHRAQrJart7c5tHpG+84M61BcNOAYrsezX
cETk8zm25/hVF73U2fTpa9n9BH3PJo2OBrQBGgRXt+r+WaTphwqlJ2oOzLlx6v/dny/yz31NgKay
xhJ4oUXS6wXqDf7TQrh0gvrKkMIilbvwslO/Q73bL3IjUXouE16sKwB13XDBk/fs9sQbl4PKIw9t
O390O781tknMPQ2dTIlUrPPOyyx07k4NAsgH4rUqi3pVKkyoGiwGoi+S+N+/mh8n6Sv3/QssCc4x
7iOCYl1M0IHVus/i4D65Yt3T0HTZh+idWyE1GIX+2Du79ElhbUGa0+MkSQKQkh+zAnigTxD8g/1U
nMVaBkeh8n5+KsXH1EebcYzKBVxFwYZVMyQHoIwXB/kR9sDy4XETIbEqPB5jz7j87nHEJGunwH0k
smuceX4OTpv9RpzvWsEyLzvVMcQLDx0xzkXrx+ep5h3YJQ/bnyD7o4M6V4ynR8kkvILpWhqbhnO6
5aFIIX/6LlqkQ86J0hDt4+a/J9vgkJMDfJSQ19qb2yQYEDUeTEhY83Y3N7gPePD+5bFboNiiR9tY
SZA8/EEvxgbs1b+dMCLvQ9h3VzmnrzaMywDo6ZxLsS53DZIO1nYH+naxy7ks5nGWAqsYDW6BbpM4
CsuFgq4/FBVW6lZGYW/C3lDIVdG+QNquDPF/N41mBqkqT9Jlrc/qS78peHgYfNUkjA+YqTQrsScI
JZBvwal/Q6JHjcl2xgB0sdTsctazrTpAyR7qwBOFNXfwuG+LsCavD5VIqRqTLUdBxQbVujrjtPyi
6T8pmvmslEjDWzJcvgju48kTvXtvCiEOowUlMIJ7SJdQ2rP12HRRCHtt56MBznF3HK3Z1QTysfsI
mdBroFDXaYGgpLux9OnaB2eU2+TQ0gAHS1XTltNOhytJQw1L93oTmPBtfovWk2bVNqLo0DeaRXBg
6NA6is+2BhHTKwWNaVXaoMu2eOjzUY1Z5ucc0c59XYKKpCDRyGxhOBwB3aFlrQ0xRAgIfs/gcV6P
SIShAY5chfpRvWQLVpQocUl+DJobTJE74NxQRcEMJaQYgmpbL/PdYB6e/Yw+BjsG9jDpUvb490AD
4HIcDvSGdX9Ancr7d4OP0tEHu7CNptnDm6YaQa86IKKlkvzqf30oyAXCyNX8D0rt8ynQErs8G+9b
tBT908zCgoC3R1lSR55WYj5BgL7UuAgQQn26qQjABumhFdzMndzvKSgxTZicXGdeco6d5Yd0lY3I
zMetljOCx0Mk8Fom1OOwH2YLX4IGh7CL1xb6mddgjMR/iZjs7bH+ZfdEtyGVaMIZa7370V+xh+zo
Ix2UkqH5dOeRlko4TDGnEB5QpddP5Gq5FZusjrOVFWmUXsdqaFqOif866e8w6gMbFLK62zqaUyDm
ZrKS6dGvwNbxoVNnU0HUsM58jpDDiGo9BXFqxeoLGfXE/la7a/SPEg9cGoPQGTFpyggnS6ga9IUB
ko7Rm5NnrdnwA9hbVF6sNtSDjkS2Pb9t1YPb4TPhB2u+p0ZbWFN67aSWW8ctqT35KfPQucdTVwmG
XLhPqDnTqiVqr9LxqEQ9YQKxhcnv7U10gXFAsrAguizkgieIfdAj+5kRzpt4jCT+o03xuXNKThMc
Zr95isj+aRdPXHtMlMYRsL+tB9hE89WcdwMHCqr4kUbC0CZhCh591XNlbmk3VROj7p7CJG2R8Vun
LCyPlwbiT0MMFmsYdmbflL7bjaIk+7l3BQHB2LeVReDuIetbU91bFzGij0MXxbdea9tiyzx3tMeA
2ZKGftO0nd9JshyNa/+Pa+wcGTZj+GiwzoCqVr9rdT2ZwYZRGiQUF9ps64ZpgTb0x3vKnoAk39Vt
mk6JDItsiYTaXQy7AbEYtorIfcgwx2GSwFiO+ZFHrtI6VTlAlOI0xYwqhP/hLlEIlXhXu6CfUTvX
8OqMmFw1qOoq3MwadYiFtAM++qb/8P0HcjzrhXQ7FgYCL+EDy28Md031aBk90rTDPi7X0uV+TE1E
Bk94gHU5M3upHUyXjdERwyXA8um5ATPtc0lEzPzWsUhX50bXhxSjEfURfD3qL9yZnhK2fiWrhodw
ddwPKyaapmQhYRx7b6sPD8ntmH214ofdDmBigcmOVTimfogQu8EbAJeX2WX7HYhBf3CfDuBj1896
DmW4EVZoohOQ+yy517z9DMaAuMhebx11ANoN/Kg6fkYbF1nt9gGcis6ePjrUc0REOGbO7GXXBNld
73FybUWJRGP+wWZ8hdvHeDqd5Ct2WoaYCc8Ve4tDKUmRwc7BorMnNtGcvghzolHb43zE/lP3DxMw
F4NK6Oq49P9tUCIMjlhG1Mxu438nbTxJz5lYtde4KhBBFf+97b3RJ+mfIgmxj5T86/v0UY2FiPH7
bCnfEYvOrVw1SWOkJhCFPE0/KbIJ5WtLiRwNZxIUikOC8AkdQjECakksRbv8/dAHzxcrh1aGBJXr
xaPD9RJpDRN/FWLN2W1GezJi+iKo0O5guddvvVyW16gSDYHNdCDNSMEW+eCg5BcFn7/EEgksB4tK
fssOlISt30zrBUaazoqalGneJIAYHYcpintrdtLSiYmI5TfMELemf9jOB7XuS3WUTLumxnjF8YRk
53p+/nrlwDhwogB9QjHWiV0ObDWmJbaMsJRHO5e+m4eEpB7XgMca2qg3RGA1gPor1aFRManmGmNn
tOcUwgsiYMhesuWaw69/L7r9URp8+vuOEdftxavaop5kZ4rZQIMiRvPBuhBgwfmjU601snCzO8q/
jMNa11bXFv/+DTiyYy+7OZwdFj2tltUrd3zYCPx6zbxBkzEVTLltCDeAn/faHP2RfxcIN7DQNTRE
vjq9V/snJHptlkQmUGgOg5TzcE1lsD2laGfq4Sg6rFlg6jp5kyS4t3s7B694TKa6hLccSnTpQttP
3NathUYU5aaWwZm6QOmiISzdbW6YAlsIuMDRjSlMNcbZoQ4OdlRTzPG1gYn6Y6ElOM9wigyQxQ9Y
8sjkmwSqGeI+Ya3otcevpB9MH3dkWS4h8BcrOKzzPQDFMhxjHkvY1UUPuSAp5J88lsf45HBqK2ej
UYkaFzj07yUrBckiB5DlJvY+WWZqTothBKvaQT+QySXxBjL3/TVAIR8ETegdlne3aJuxWp0NTZ+k
d2OrSZQGyJUxWCkFW19SsAEoTk+4q8YSqtuFJJmiSJsWd+zIMb0vxzuMdhHQkMBWaotTvb6Ed5z8
iyJEA+dSOgaP9PYobPNHB5A29d+QqVKmTj8izMLNaikbYPzHMNk+X6Jz3D07WTk0s2e6FytQT9fX
ZudauV2m95mU1U9zoP0Hi/KtmLu71cVCw9vZPjRbdAw5T57DOlWumJq/LilUgEFmX1StqNsq0X3D
onJS877h3csnbhoJsx6FfNYPL3tkwR8S/oRbq3MpCmUafRnSqPuafrggzQAZ8DOUXEfHf9WddaB5
2jXF3FJ+Dy+YC5oiSqtJb2732eY3InfvI/Y2DMm13gfjIV8pwPpX0gAN0SSJy0SxrEb1hPFriHvM
ZtLhMQARmOiQ3bynBhrsE9jG5WUVuqUqJL+xo8EGJoURc7+bpdVeRDnFdGh4kZWo4p0/uhcwCtIF
RppF0pRmpFiPLlHh2Lr6hs4csipngVg7FxQKsWHv7v7IlMWZG0FqFqNea+nNOH538XM+zAsDdBbb
aDlSGsGSvJcRVVGHi4+za5zkOROVK9XiwAwhwL0wuzTTRwNKo6K2pE9X898hFjjz5dQjMegfYNlb
T6C3p/QFF4zm5ib9lcxuC7mpYH1cJY3Bn3Pzv0I56OFsPdl0UrfqbzV10uNnORsZ75McKZk9FkFj
8Xm0SdNvlIoCBd5h+nOX4THWbtLjyCDTu3ZZZrwQ0sq25TilTlvSVNGWHISBtVPKkOj6OAigOrF0
rpBFrxMwTtNag1ke9UP9fc5eZrV4XaswByOqsLRt/20mIkgInejRRCJP7O2iVXDvwlRuUvfneez9
LVOGsER2NmkkoHL17pVIa+wJRYO0i8stABlkSCw5DmejKqxz6jFrBpQvJ0ztRgw2Etc3x4QlK4ER
QIUsbMHYcsJMYhfh7mN6ZHXQygSPEJaT8fehWRpSee70UdjRBaLR+VYZ033KFUbDJcielBp/K7kY
9O+pvcT7iHXM3LiGSPCNzpiOGGvgIek+ppGQbz9SPlNfJhEn+txKZpdTBOqPOEExG3D/TfpIvz0v
O6eyt9monzuqmzDnQSR8LroTMc2R9AANL70VnhBA7bRw9jvLdlXizbuD8hELkNteoAcIXVGcTkfb
Eu5Mmj7TjdQac9xsNy/d2aPHaqczV4oc77BKiz3BnpT9g+cmYD15lrB8wHaPp9Kdl9cZEGxImX2g
jRvwe60EVr7h82EcfGsMuwO46rnPYeSATYXMPNACQOZzSH0nrm7jQQU07oxx5dNy9Pesbp3aACqx
uA6HYG1E4yG83yNJ3hV8YL+wgRmiyc4QPnoeQQtQcNKjQ9datfoIGsPACU0mYrUOYYELJPYMz/5m
5nv//xTK2n8AoeQxL+I94fozzymp8bvWfkMlF0Ga9nbNzzCMKW88Sw/FQazz+/Sb89TGUaKFzuxC
WZ3EyvrcLZKew4nBS+idUfUxOtxz7Q2cHsVvJ/vxy3efEIK3S/pLGB/226AeV9TnkwN3pC5CcJqG
+LvrTeBXz6G7Un+JcuV1n33Nn3rDVLVQiEhRW0S5IxeNFYzjPQ3av3qQqaVtlIE/j+6RdNUTKyeG
TZ79EcXtO02TtRtqdKG38DIkWg68tttyZ6UVNof3iVsYzwM93zTbUZ0OnuZLoHIrcxVD1/eQtkXm
Z+DiZ79gizVjmTUrHIKE967iWuPBX4Lr4l8roen+3BXRP+penTgQG14ZsbSKvEz68fijdEdK1RnE
PR/7nZ9ecTaIjXYfQMb5GbBK1sPph4z+1QdfYWMtBkljKF4nMI1jnWOTJ9tf3vshZw/9/PiNOxm/
EPqi5bi1ez220VYjmq4xidzghvsfoF3Eker9Lw5d87xkZvIfx9byNb3ah8XRE2l2+cCgxpidtY6l
SIofiizSg3T/t8vPpuA1LZ/FMvMO0N+jn2Py/LoMomSQm/YNjfSEGwPd8HER/bvJNw++cnn2kTX2
eG+r80NBD8DVMmAIbCVjf+1NSoK5iktP9zv8WDHZC87KMTGjYbwPaB2o6Cr8X6srsQZD1Vprxm96
2ANvjMqzKgpaBSneMIdr2KJB//ESQoE9uMAI3ZCsvi5TmEogwAsE4pa0a9d4FRKF2SKYXEwwwCoK
qqkhnR9ZaNTSMarCYrmhC2dp5sJO+/gJR/JXEGi174oZMpFHFKY8vSgkoXgdf13Cui/NIpne514N
ei02xbBv/ehiRKUyCJkKr2PBYM+Vc+2b/z2Gasiw+CvZsj+d0mvJQ8g+suuQDg/BLcyfa46ttAaF
zeQwIs2BnF60iX+2PZM1P1pddjtH8rTCDGNJZNt6bBY9WyXS1yoK6DRY8TnzSkIu1gGsPA/0IROO
WNkIYz5L9u9MT6jdrJdUTiaWZ+GbD+qOM8aU9dHzH7kIB37Vp9amwfWqpWRGkgf+qst234JsEJVN
YJ9CSS/346e3EdJHDA9g16qgyCccx+TVIbPCB8kfScNzGnVWmM2PhwQnnzUUXeFqyJDjOS6icJ//
g903UKa1QGiZkRCtkCXPBTU/gvgTsYL4i8hC9yyvVRVXB1MiAM8iDOl4MmA5OxQ3N2LT7snnWebn
q0bKw7Ci9AT2nI0zSkWaU45MTptFhCOM+isSplOuHi4F57QMZOIUyzAe2AyVOyl4csPSTX3tYwEN
FdfmFJ0RzdTvdJzZtfLpIJ6HBZxYzKCGlBLGfpTCzR5TohhhrK06uKxhYd68+av/MydQFvMg9hs4
4N0pNxa7wz1dAI3JcDZBX3V77Nwkr7SWtFXAPJ0XfQvr6cIpvOU4m4kVYGoruqnY5nayHnj6a5ue
UxYaP6zoPWcVyDT9/1obW8qtGwZOneeFg8SpAcBPxYpS+CkiCjryibzRos9G1S+SQUvDIVty1BrY
e4q76bUVw2ogQMm5SXgujjSWXks7TJX/t5ld88ryl6ydr+9cwur9biJwe4XXC+zJsMCq2pLUdkzw
USpLfXMKulc6F/i0VzHljcunFYvMjKB5NPRJAHFVtRHGuT3hHh4y8ouQ8WYBXjibXnPYIf/90w4y
kyeyZRlBf8Bpo71p4T3WOXmviCZhnTiWIpxseaUJhTX3FhOub468Gw90vgiDgh9a2VbQtMTtMZJl
k6UL/0oLv3ubb6yXR+rGT6uoG+/Um+H1dFBMaDus2eQbY4Gb/b9xYybEsTtK1qf2/3g5lBfxXOIW
NLotnR3cGWbvt0FreYavMitTYzmZ6twkIDcwWFPJgduWLive12jZHazzFjqDgVpTTKvl3j8zxiEO
Ps45Y+IqbCoK2XlFzJZP68kaxza4xixE3BECx4Ae1ve6s+gFxV1RT/zNtvTLqMM18biO8zq6Oy4+
TPNB6k4Pt4x1opSh8sLs508MgwVhm1wiFNNCySrQf0RLqFwwxMuRdrEBL/wbuJCyeEC5YBkvye89
7EAkFCMu/KgUdbiFovDQnL4AkL9HtiPUv1WUT+g+N4By4mZPpR5XXOdkeNjlvkQhWzDwViCINAp8
zkVQ5nKuLpNmW24shdUctdMMz02GJ1OtGAtxFCFN3t1oieYLcB1xhp43hpalOanS8Q1P3yJnutIf
II8p7Q1UBV75LwoD285xquMIlvn0f0MC3BOi9Y9nhDh4WWGVjZieMoylqnfYVBA4/6Mh5XGN4Ka8
a/u0kp6qbItm7PSmytZXzSy4qX9uhXqPM2qqPtYpsMUcrUvY+6WkTPMJ2hUuTEVgHunbfuP6Lij6
07mBQzB5orBtMrtsLKQI9/aqsrf4I+8GmVsT6pvlCjsRWkGv6dZmTAVdQUlg4PddgtpGtOxPww/S
NXP5e/j1LzdpJOYq7eV6/HuXp+ZBolxTTiDHNFoltN8oPyhKgoHgrKkF5ADLE+UO9pB16QSKqQhM
NxesKVp9nw9uo+GrwehUlIT2zGfLMDWj//+BtaWzPYZ3QssyMoEI6hyYqLpkYRPddS7HOYd6FxR+
+J61J2Rp7E5tsrB437XISLGK7m9qU5KwFX8WNhrdnq7zOCNlYspqYCs1X/JLzh19v+FXuNv0qAEP
z5VzTOxRh3yCAlZGLn7NTF/lbGjk9nwzDmBUxdkgWqsxBcSXTkGHuAx3eKbvm4WwlW+CzdFwdQGF
m5eUotNHJZDARvDKMaZxZNFMymalFuTcrbZ+Q8oeyU2H5FW3W+PWJ4OZpjFE6y/n+Ao11f32qjxI
1NTulJcFmDlU34r8uSEHhxhrUj16PkzU7nVi6TU/M8k0hsLfLrIaJEeQLW8SW20g4GVMMrs01rza
x5+xRMd5iGHmnPbN6OKp7s2omIZK1txw57MWmBFu6KFaExVKlbo082EVM1n2bpFgFzKoF/KwPhFN
fU60gbCfDYYXUzKSp1ttsmZ+WLV87c3eDO596bf3zWuka7YMqhta5i6EaNbwpqRiEzF0yhj5K+Yj
BqGupkF2q6EpadxinLAVxWV+9ljX94jKsdMTKR9pV7uPr8n7W2/7kzZqjXoKhAmu3Cnr0VhMDSrN
P5oNfkJ9/9+NhrnyMox3lPjDhQkuwo/7cf23iPCclI2cRE7WvL0xqfINVlz4tR4HxLaMPyXfsVyo
8OF2d0CXoqyiuHy+YD36q9hJ65qejUDp2Z7dfepMEvSi7vUJt4WJZdLVLHop1+xhrinDF/rZgOPx
dQsTbughBKBgyciHAmnfC6KgBpQNio5VlLYjuglL1fSGhCBZdReqF9vF521jCUDUuEiVFF/JAQJE
jnFPM8yfx0vM+41aLlZ+DndTmKZk7JMbr0uU8+/5HcFCSc07lspljqKhzQ0/TgJT7fLrEHjtjSBp
sNEsQv41xkpbAXgEpMO1omSbZFATGZG5cswu74NLu/AVCWSYT9TcgZjO8GjRBEB2QVOStQMg7K2b
WmfOw5F1fdTjVJiqU1cH0kPyBfLV8qEpFUcMsxXs36NpL8a66KQ50xtM68CXqygcBjIiejs+ONQu
bkFrviJRPdJo00JqjXViErC3utWU+1gOYSXua9C+TEtMRWXps7dQQ4WvvH+YK5InLBCrmE+2Imn5
cmjA+K3df4Uh9hD9nlliiiI55B6o1RhUV/ajBNbaUJ34hv2IXemsT/9ovDmhgJMwKIDrfzys/ZxV
PaMAM7PQIHHp2om40PCH1WzoiKc+F49YlKEn92sG3ClNploBRz0v01HQ4yYFX3mE9wcrq+147JJ5
7kW26d3vvHcTwg0lKDnwbpuY7oE5VCvh6zxHWbcwtcW/sAS9whUrDQmUpA75Azu5DSYpj7ulVgM+
vYPlcs4AYrzfmx4YYcpUY500ombEhirJd+XCS0pNKA27qQsZqHqynqGO4o4wK0nIr89HNvwhXj+7
b4l0EXU6U6Qld1zoYUtvMRbFlghmSVzeIcKvWNp2r/HY/OQaK39AS/shJ89j6CdyPus/DIm1cl9b
OVskpNZy1KF1EoWYv3TcBCdbNKvCbolh1z/WybjbwQl6QgakJX2dbq+IIgU/JK19E9xq2VkRrX4n
ozMOkj1UylJgGX+I6gWT4ZoGmOtyRMr2HfePYM2BaCyxa47LUypeq3FrFFB8kmHIi+uc6PlxYXCp
icDAmjVzVGHUraJeojYfjYnLb2CmcVotxUxkTlrVwz+E6/O9glCA7TWIopxm5rKNOwiKEGLi/O8R
PO5gu6kuy/L43KElaB749i8c8Ty7HuOUaDTzjodRznjQzY3csLBl2nhqiIRb+YfbxPY/EyplRQej
96uP5WyfI8B/vNNEgxr2VTpeoGs5mVOOSchcPd3qhybIWCMprIUUOsQCIv4GmOj/3m9lHor7BzjA
TqPfweNFnqSop6vrK/Q9uzlN7KTIZra1LPcDilkRE6mQtlWfONeDODJ8Cdhlu/gPjQ4FZaUVI9YB
HQ9GZtl2Q21ZPNBl/d9vpcPFs6jXnhPxnuz0bISMyXT+DSosaGzMazEuwch/6pPgXACa26VyFz+n
JxQUR7nHHaSJx1Xw0dp9TrYtwxSLqKt1JVp0gQn51lwnui92WzJT9kfyhc3YHRxz2XDjLcisDmAO
9FWLVR2yzoqZMwu1yb5WYGOfrtWl7PxujOTZBq/VWE52Uc6v4luDQhK5hHaPm/Vilv1RJRgqNgD/
50kPrmHuMzO7Nz7AIEkyiCWHj3pPV7//3XlEXyn00nADLY+jQpuWzCVgKfVsCKWNhM0bDDCAogP+
z5huFI4AZoC6ugsgYOEWkSNVyZgPTcJg6tZTn+mrDWnIPepZBqzvFGWzbBEt4tR/JWBWwde03tGA
zgL/ezULiC/24pv1x8BCrxZTdwtiNWP/GhFhzkD6mLLGp4TN/AwhrDIIpEaJ5WsANYULCLObsN8u
uDZ8jP2ph1rwbkUwlr4S1j9S7RMQEkkRSltxP4ryWlf/M/I/5KeisXQNdXvBasfUZV7yAqiCPqBO
URU+HKSs43dx9jZ7Etedlge7Skbh6BwxxobubvnecuYsksF0R1xqS+hHBDedxJCOfwIym9UsvtJY
72JSgjncl6W8GqxTQu9Rp6EVlHzfZMKyPKxJ3tZPmdsKAewvotYP/jcIJkvRBBxEJRqZK/Dw76+w
af1Q0NAbAsxWMObMfO93B9KlHF1AOobiuaSv4u7haiB+URlArq3CimGI9PSpeszhmo+sUxB4U/FX
Rw9FRRDdaBwxE3SubYBDBCAs2ARtVRCZ7aIDx+XhKICz6/pZmrbNjrxZVz8ddJ5zaOMLqfjHlLTK
yYKBCXLvE3aI28VmDlF17mCbGzBw9m5nwwtYMaZhJ3JUGlA7y60oU32XtBtrPRuM2o9pAULP5/CP
WBnaiP4pD3WWHOyna0GhQyixh4Y6XcF5LZ6iURX2CZjVOhONqCDikzws4JkxeqR7w9zzx6FfCoWB
3gOip3YL+PgBgXAVSHpxV2Gmk/tx/aIBoAQjxLpKDrXcKVsToj3WG+vGgWeXA+qO/uhvUlPZrijb
eCWwciaLemQvFxwzdIysiVbsSssLxHL5aQHINiGYV8BU/bE/O2RAcUAxhgRGW+U7EbXdkHa8fYKW
06g7WZk2eINUo8vtHqNU+CY7cjZrY2Y+uCWxE05v31Hh6shkUWfo2et554RkxvGqyeUO5isq5Z/1
IASL6c6HKg1PsuzMY8cxfN7+y5sMi+JGc8ODD2uXD2qhPwrfYLlv3bJOAA+4sGxldNUqST00r4dQ
wRLoLs9HKdPsO4rcxs1mMREbL/r9dJgoPYssb7D7gXZ9gKz2mqOTM1jhdhI4HD7nbXjoUoF6O+FH
RX9DKH9L34Ynn3jGPvoLQlHrT9kNjOgpWzSPEhEk1Q7br83b5JmP4ka0B0tY0KKx+eoBGibxZBLS
XvDupUSxD5pbAfLcxcEmQ/PQcn36aq9uvmScLKgiAV4cQ38ecnbyNjfbWnJ/Ox2B6QQ9mqZNxsaP
fvHNxqXYoN/hmmMIOuhD/XIj/4tJawQuKRRKPHDKG+8CEy4YvOHdbCQpS7jSUBlr6b+ME4pCeTQI
E8uVT8FvVmiKeEhh0ayt1jJn5H9iWagYrSAMD+1y6rBWLf7yWaMYmKdKln3dBUodMiqcRyBV8c4e
pl9oVrrVENAN0bZZv5TlBXg1qYMteRabrSuZahOOmj8F6LThnFg4EkYMYRzmK5eZWEeRDs4k2hWc
PU/xDU52+sO54R43FzKvIrjB/yjsJUG1xktJ2iXlHTTGbx3XDSgFmDSOZ8bomzA9d2qR4vtkuBjB
MhJT8lTYiQqhS8M0hb0njmMO0rRenjqhSI9g5+xSeVpI61EZkNwrKrjCiIbYx1HLyLRo0h3UFMts
vAvNOXWLJPswqjbSdjm1fhgAAq8Ec29PptcSB+ZN5FyWrfEWmSILQYhufpi157cwgGD7GEuYzGjm
mMS1v4jq4ntEg3JB5DAsepBu7p1QhZQDqH0GRBw4ZzK0tr9P+CbNanwdySAKCBSvp658V2kxz+nG
Jz2mf3WPhm7fSW6FT7yqEJ7kZp41ZwqzHboNCSLFDxlPq766RjwsvAgh3HtsB5ZlDIQ/RKRraWl+
6K2iXpNzLTYzq5aTIzNU3CjH1am8GMxhdJBqihuU+9nBMDmsGTfmZtOUMlOOJSj1Dn9s+wGZCAMS
GkDYIHZLcCAzh7Vk4wwdXOVdWhZdrD4Rc1ariMhaat3v7llN+xipQzy72ytvBIb/l4AVxMjSLeTq
VBX/gBPfRZqrWihq53fCxpw5ptFXTMWIMmrt1IJYXYLIKdSVuB7lx7Mrxnv7hbd9DSqo/GOG66Iw
ZW5x6n2yNnFRAcaRp7ULzy7nX0qKIldCG2t0zUiEzTy5PTFs/IAR0dV+//oC9N6ENkaI6PiwK/cA
9EETXKnQmL436GbVXB6ZfbhZFrut/kNVOI8y+yF3LxvPgY8jX1BWfns41Ph5nzS2CcFcuGOXYJVL
uvn42M7x7Ulv3EkCqw+Tfi9VibsLzJHAPcoT3bFznnzbQJrEWaA+gWkdqiXtVDMhE1BOOPakR75h
CAdXbvgC/P36QPcVgpcbuMoUOsUBUdDfsyaiSmJgixSzgBQU1vNcNkJkVNcIeb4EwE4e/TNqMLzd
LpMSdrlAcDwv8QgSjkPGTazBlGhxRttSGmd8UqDRaE1xo7YgkDm9cqUwQvLvA3kQCggeCXdgmLbT
6JGrbFOlT2jHjP0EVrt0wJv+8lnxcKuqdL/HA7FDZOoSNWCAnV39XQOJf1y8x0eUnZ0H4wsK1rMV
k8FzK01ldMUyZo76utNFbzIp3h4Tr6Zr0qTvLd9vdB8OVVtKBIwNaDEwffolYrSw+1zZ8DiiZlkX
YTcEa6F3JVVFkpg4HDX8p7ecUtWjd9VGkPjgwTCUdLA+QbQVV1CkbXcF1TSb/jXtDMqDRCofzpbF
VRD0Onfr/ycKVTUUjTWJG+NhrddwZKB0tAd6Vm09E3u9+jU8LhviY7Q4YGmQYc243U5S8to0/1A4
ppBubuB8o65FwdIsZriHnMn5TfmSa+6mgxw4CccduYbai2+p99FMcfin1ij5Kh/x/BKD0mXZT1dM
Jm9o3pflEW9oqzT0ijOWoAA1W7ZWOytj4cRBPuGrnx6hJtdGR6X2G8vVWqkn900mFoiQ6UlH4k8x
QrIt2A/PiqwFUwxRRny4D9edsvsraND9agU5Vzc3JuvdY6YVMo1xQbYaTv99jdvrA4rnxgWkEkhw
pKf7S5HCa+Eof3Sb3Ai2qFUtWVhKKv3DqnVXQqsOG3WqLw5okn35EE9EIiXo47H2cpsNNdY5peEV
RaR7GPxf8CJpqRVUILxQB94YIoilGDfbVmyHeN0/UdlEtFp2cfyDxhts2pmXhJa28TOJiVtmQUFt
GlvMqFxCfbR3yDbKkOXRShryow0AN4ahBGMCzl5Ws+yH+5JIHvNmRgc9g+AdPLfwzNo2KWlv/zVN
FUAxOO/qlQB6H8v4WFDpXU03xwez7JWbg3YCRtCZlK9ZZZqE784msOZbDNKM8U69mAEos6dv+iwV
uZtDfe1EMmfpoAxq7ZcCyHOyfwKIwQZNkgnaIQOyt/2Akmsljt7RLCllZoNCT3ciHYZAadKdgcHO
JA73JZR/fx1vF+OyUksaZQ9o4B3fLrhNz5/9laDELOMHM+rcgJiqL5Qd/K5oLcarfcXXyNRNWqMI
UHaYH/4VCJz81YE3a+ANFSN8/LhpW62OfZPsYH+U95JDZvg3C28a1VbmAFr9IokQpOowYM2ZWYda
D6jt4YRPw7USz6qyM0VyaTcUpRH7Wm+9RE8yi/N1bGaplwntw/jYxoSuYEryOgfFZaNsF3yJ2kK5
R+cofak66LYqVtFgIDLT71am9mhXifcLgbHQBiEsYqBPpX/RIRUoqqiqYPKpoiy7B93mZKyBHhpj
hjsdupS/kJq2sn1a1GLFTtfJwrsqhfGBDbMOA8ZT2j/HYo1cD1a9XSO5rIwsnDARqgZ8dQa10S6I
YTTa+0PY29cq028kJ8j28UlLoSTqfeejw9wNKAmrU0On6IROBDxDOGKldGzWxi+zH4gFUQJl4GT6
96HjIY1Shr5sGdVuVry1iWZkSJq+3fn1xUUx5tkwimxJH17OQojL3evC5nPWCquWDF2rEyV8v/TK
CNlhK/gP1yImChtn69Vs3asDiAR3cB2AIKX0ZOgcefEbwyrHKYy9JJChH1PPLe9Ou4JVUsLXhSgV
7PQ9mg2LPMf+EDw/YbiqHECClFfjuxqaz7GKihO0LnCYOE6Q1/Ac2wGSalChaghb3eK4gKnlBFnZ
RFTptZTROdNApKBP0cFYpZCTUsUtfOz2nIpa6A2th8aYuoj7qFRX5GAtRJayTCvWkdvcRmKjpIso
BmFu287MYWrzEGGVkNP7mvQBCMAxadPsTBSvt8B4BKcsXaEzb+7Fn5TzaDv3iwRWY8+gu3m/VRsa
gJD9lwd6QGw4wcuo/S0VTR2VYPLI71VmWR5oGwyPleIANFtzn9i7+LLj7iVZc4OMlodK5OlH3Y0V
O/M+TkYdKiVyICsbZTxlTSNIx5pSQpUiDimbPdBLFtHMXnwHqbbZK98sSsENQCWKT1m5jXrCI1vz
L5xHY+gLr2cuER4Irgna1YWPOe6M5yT4gnGksrAZ4y7KovDN2ZDpYODJLTtG3Nu485r1zNIq3PP/
Q3c/IJx/g+ZJnLIzwKRKly6c/pg5CnE+fFtaBdPx3MYYcj5MBWOG4NBu1pPyaDS0LeXhnWq+dThJ
+Ngl+OSmy7IG3EkDFlrA+y2e6tXf1VtT9cdTwP2l/jb7azVIWhZdb1qE75Esi9G2Zqb+DrChe3MW
WEXlTe8y0Om5nGTeSKeqP4/plfeTmWCqUvlb68cktWhNeqMjL1i3UDr59WKF8avltXZ58tQoeHjn
7hW+LYhmgcHnMi+OydNsvb+JP8AUf7JjH6WHHgnbJAhmLpsLgIm4Z4bPGLnTtQ9C4OTenzZiJwdx
AHDhZtVtJy/h+SOrrxSTU6+Htc+punnm9ud32UZIsXycSDhHqhUi4z2P5Pp9Ffrb5U7RN2UcUC5Z
CuuS+KFlUzehY744sPWiPPOF5WpnYPPAQlT32kcAqmYhVKaJPYUBnKqCwBN2T0/MQPT4YmmG7MEz
Ky317u0Y4tUY8YBYzIedbPnChnpPY0QpvcxnWxkNWAiXByqruWjJi7T5HGOaEuF51CWegUV2mTUv
/XouSU6as8cGmBppqNdjLFUWZzuqfh/R6BF45xWRRW3hsg51KQRHGVytcRyAjly7nPdazgO0S0AT
dThNsqsVJ7/6B9zBFZZoli3eb9qSbcM2xLsSxBe4pDqnPso4Zf9lbUnlXh9LiQ6abuuEhjZUI4Ve
zkjXUafnn1NbZU0AHS+TPHNUJvkUakNgHxk23tJKTrJy8hSjhiKE66jf63bpd6H/4BOwT7k2jQOK
+h0k+ONlsRJYqTBXekUXN6GAyDWlChLXbN+tjbGz6zToVWCpm+e1n5wiuTIgBLPtCcZbZrMFajDq
OjV0NV2amYJP8nosk69zttyfRN4wm7slA2ifh9tV0yspv6t+V8vto0EBNuJrz2QGFFOwrEw3Ku2C
fBNAI+IUis4wA3doywuC3N79B0JhosS/Nvc6sVleV+FJtQsyq6U+LjNSk+MswSzcflMCfLSu29q0
JQwsnYPTUyhhw6YD8OWidCktOBgTMjSai7SwUbLGjcY+J1hRuF771zYTHthkcmeHQPI/rY7MsyXG
+VynZYeyAT+pW6I8EV6pPtli7mCTt4bPexNlN4S2NgvlYTzQrneoCLrC0PEW9dQkBk/UDwRHbDzQ
7XznRUFbyDc8t0w5/KH4ybbmZj6TdKTdpB6HEaBVXL3baP8fqHeRjMHODxZI013sNLJCZMIkYDSX
3jnGfpHJ6XaXwKWu16pKWFyDENMFIpFbhqLPmbNkGYTQUMe//THyx0O532R2m3VggK7OMpLe3C2N
LtrOqrzwTIimOiOg9P928l46T8NUrskHOzPmP7rCqiTgICi+Ts/HyDEmyFkAhFM1Y9AZZ+ahbKOH
/Onz/o2NVAeOQQvaSiaFr9XzwZvyE/cdtCax3beqB2RfMP09UBALkT0KDWPn3wcJ6eKXpWnSZeT5
lygPMnoLlonVLTHG6g5qHzs8d6zlvgsqwhTw38fVL4IpgnF6YoaRfsGGON6EcKsfb4bWhIF+yrIv
+wSJAWuUE+pesWDLQEOy9FVGQY6YbH2UAPBEQKsHqDvda5b2YCO1v6umCYBCAFYrrjDWu4GR4ieE
rnD1uEi7mx5oRnNqKpIkRrLTtkZRPBcOGKr6jrysJ694mHVnu65kBriTS1RMmG8eQmDzCakOvYcm
/6PBX9glBp/MWrCVGPTFmNbgGO6xP6MWmmh0hyzYodmAKAMO7Ah2Y64IHR6Kj6U7/8T2F5G4axD2
BVifabVk5MWUAHveY27YCkgvaN1j48YdfElpG2tAzZKm+25Ymmzi0cDwkmfNmtgQyuFy1KlRhYO+
gM0ZWOFTAJVMIoihjzlzkQju5itas0H+ZyDuwqJgIq1+3kuzI0VAV0Xgoz4naie+88XfFw72BHcp
W9TVBJbEoAZDwEcdFqQew1PXznsBN6F2/SLJbO+fEtMWw26STNbtwkx2Pl7RMdXsRUnMz7bFYEO2
BKyAjvaHokkxh9eIdRDhsNcHghMl2E27wO2lfSpZJUEp8RswcV35dvGYHjPBGE8++2gKZ77n2NHU
QfRu4fupHmhLxeeW7Slp1/zBMek7/Xh0CJMc3tjdgMgUuNeq7zudg1qK5kw12QLGX8rZ29bBg0bW
GbDzF7Vg8UqRS4QWMDtD7ooxD+jlvmCz99jIFpu9d/ewMdQ4bzB4j8622rgSTdG0x1gsG9deHh9+
jOBI5uVZO6rE7kRH0AoFjnYXu1ZBIb897lh4klfssXaQ7DiV4Ln8TStTVnfSkIjlKzOHJANJbti3
SIqzc5/llrmNci67cpm5DSk6JXqIJB2EHig6LXPBmI4YT+1Fl4s3GGdBZX46vKFdzR5CQao5EBib
lH+d2iuJVJazpE1+EEEUP07RFWXFk2lB5Yz3eDlGaCm7iYkGPl+/9Mr19hUmPfyD8zQNRuewDyNL
Sd74Zv7CeesxjkbBr17EeTJRhm0eRLBLECvwrFXKTWnQSWWmX1h7zFNqeNC359opRCGS22VhpiO3
LCLF3wOqkBjRGAboY+fFd+C4V+5+jwB2fScO16/T/9t2Hd3i/wNzB883TluJ6SADSiBvhNCJ75ce
5yLGDWYPnPWvyU4vQ/NCgttNx5btim1ud09rXJHYOiM/zjdRlPuwohOMVdl+BRsNMtjMla0EXYuH
XM9Io1dQSAP7vr4OSyFIkUaSDWI0OwGelKCBFITQJ2q6XvYxUa6G+wsIgSzM/518x0bxN/nMoqXZ
xup8UgU2aYIT6WOBTzSwvE3dna6+5xSBjyth+aiqQafHjJoJ3T+P/iAQWjSgSWglHK4ebSHJPP/L
XWLZWAqJtQUo1osk9kgnSmpxvIwkanQxHIb/hOCLcVVVG/qUtVT6/Z+VtuTCYZmFSLml3SdhIzJu
GtTnX4ZAFehGzk2jEhCNe57nMwjNu2akQ/5fuH60PTEgvCdiAxQmssmXIVlWnb3Kc4MVfcB9YuXj
7Nc5BFBjb8EEMJiljQEqnyOBNQfIYPSXsSIDukaFOEaX3DLf1keeeF/fgsLXmYEtCtsTegBL64CE
gc0TSUC8k+DXSX55DqfFqOeFOQnEZg1MW/ghihurXN+mc31IA+NeRFeUeB1W3+/k3Yx9MWMZjLzK
Y9GgU0JTjy12ReTnGAkRZtqXKSV3Wi53wLUVuIOio4IxjPoE00lIoSb4inxP/Csi7kEPYfwnZ7m3
W8dvjGsRauk/1P3zwPMzv09K2C8BN3wCU5Kb4hle3rp74CnMlJFJJnU+eSlpQGRfLuGdGqBtnhNp
31pNAhZELs2aQunzPc9hnmd/yuioWExJ4qGbqWG7kjmPnuhJFmQZNViZaaJFga5D8OZr907F4oTy
thez7zs/R58VgAUWAZB2pldmh1L081PXXLF9jL8ZkLJ8hC92c3SH5Wi5Ll9Q8UbXuwMpq+/QjnhP
GrKr3/qlJrxST1T5gHpzzB06NC7LX+mstcTlykgcrxrgurkQk3iEVQ61aP8keEPaDE5YM0BXvIKs
2IktJtDSojzdHVc+qkP45a2KBdulicYbj9ik7hLKGFkJMv6F0aq1lSUptU2wA4b1QLXHh+SrnfxN
tODfUPSPzs5cKAPwHwvEFPvhORdTdAGRLcsi4eYllIWb44tTUWxJI/ch339iQqsGsDnPdOkDDNEy
VPSPWIkU6B/GKLGSsw/7bY0hApvx5699yd9Ya6dsnDRyLH0cFivw6CIQlnLU/hTDXe2j9+mHdeTP
w8KEUeENr/lNSj5/E42f0wqP/iGa51X8choHf9jffvLGxfW+mN/EzYE6p9/qMr+cAvSAPZDnvB0E
SfAgQ7+eYgIPg8ZPCGUb4mqmUsAkVVeT3mAWTFd7qlPeuvRZGq6HqMUq7HNbOxAFcm0Y9K8J3xg0
ykeAFL84GBcSd7MrMhk1bjP6ZhAZgLmsIJyT3S3GtmouGVP16CvQmyVGQS+xjz/EppoJVsnXl2+B
PKgE1aMseyDTWVitexmZbsAphVa+NXQF1KPfwYd7/fZojuo92WwEJyMyhOvj8SCHN8i2O9YV3dGN
Qxabr8EM/Ud/84SZ8Rn3ggmxWxUBy3e2uiAU/8AzGUBk4OVxdj4SFmRF/4nznTbSLzRQn0j1G0Se
T66KKxjSJBOsku95XZgB8ZpnBLAExqApHqus2wpghgxfF2i/q4s5N8YFaDbBFweRpa1agt+MP0YR
LMi6TnTfZEGF/1zQCRD+Adzz4auZ5m8Hj/85XLLT4JMeTAkyAXgt3dhflNXcuhMqPffxrnlugDzP
TU0X4FBnF53Vx9m2jhN6CouCl5WKtNG7ixIM6wY6L3dXIOXkqzsiJsGbGg69vweZOtvhkqLLKU5Z
m9eB/ktZFfXqj9cdau2jYLlNONck013ff0m4GN//bB76k9rl0b6ADPFJaZc7pMKGgTpBr+XVD56d
y3Plghu+EkLXQ9jDidFRPwS/GaLmVHeMa53hu77AAJqr82q6AeUOYm2tcZ5nswKcjdl0S2AeiHkH
f6Euli9ZjGsCTF3Ln+LZtFpT3nhciQ2HicejcHjfXcFz32Dlxak2FTTytGCHIGrmVk0pA0K9HkuV
INOL+4/1j5U3dXCQcd7JAFOc2Tp3kmnX3N3+xjqJ5bdxcWg75iHH2AmfrKQz9nmJC95hhLNmBCrH
VB9CepVqydRB5cipmn4Lvks4rgOBvdFvSuibAkymrWkHTyprR4Q6v4M6YRC+tivCuNqW9+I+o+7B
oK5JVfrD8gswapWe07saqREvKiATbY6dVKw0fGOYWeqEYitoPffbqw7BeSZfdXoXDo9Zu8z2+HDX
O4DdU+izj241bTh3iRywg65N2qdmRFAj5RAbzN9iJS2rvfudVNl/oKXhDMWZZx0VODhH/kNwq3r1
AfUVbURFlXyIowQRFhFaAtUc9+uU/lydJHRz2yCbKGB+m89lKvVLy6QyMyi+UVJEemhAKBEeRKdJ
FJckfsPenERCR+9hNDOgz6pjuXGFKNWlz6YIV9yVXSUdZpdCApWs8t2ONW107qfiwnNXI+tbwK0D
nJXgWA3Wr2FBvi01eZQMr1+XyMeFyrJP3n1yC2hQMRdCEv3myHapj/LEROT0PopgQ4dRjxQmCsT8
KvaK+CtEB0SMVJLQQTjGh81jKepoa6mrmK4tIZlpPMkhlGCWfOIvSv1BuHKnbddkKiYHrgqaoD0F
e7f1E2cvo6FKaoYKkLa8xyd9TjsGYqADtO+2uro7WHhxrvS6xkOETb1xlryTbgn+uKBXEcfHouRF
xgDTp+44Avrz5Ifsh/l3oCsQf/qyaGjxYFCdwdyDhOz9/YBuXCSMyou2GilDARKnHyTe7oxinp8h
GtOo+WMcUYbS2B0Ro6rewTquMOBW6Xxw1f/EjmOHdORs6+wROXb8vxJugc4P8rmauj0rOJwMmYqk
YTO6/SjsWGwBBFuMr9QQJ6xhyDHDlLCypKsONdhdVunVthdEb53qd0O4kL+8nK4On02Yo4GrPvHe
pJKYcRUb+rnLisVSuuyqlw1LkLhpsiiNVRBfqWcFbdxlTLAd4dIwhQ6kLGvrEyCr/UUHafbroKm7
ThMDh23Sq4aoTKgoEnG0PAzDKoAyCQ3lrmcJSUO3WOyspRdm0FL91ZUoPn5G3xHirbuKN3MdWSmw
4oJdDTC0PB4AGNdLM95CYvRFoSJwXOeMrWdVprMhEybTkvj53RZtZUkfrR3G6wGheI/41Doilr3K
63hkMidz4WlQ2/xtSobFU7GkgPolvhurkL67C6mlWEdxjGBOQqoIC58Xo0/zBPf+cOm0udpA/4XA
ksLBls6cJWYUMb+AVjDFC178KZO0SZhnCR46imo5vULkR03nx/nv9Lk29jpUhXuwzqaBTQ72jwDW
0ewyQjeYd6ODqkq1PFFLO9oaiSCqR6QgWSq8BggmILuCf9WyecXyOld3q0gin1sD48a/Z2lDhpka
ZtijQPHdKDFqrAEEo2FDNCpdcNEHGsOdVPuhtwpFERSbqCoRX2g4n/D+O8Bkfm1qEtM0kJY1mX0K
6CakuLmfXJXGHyfTFpxXbaIWdXjEXgik+DjOk3CPDTbnuXuBMWKxNYwSQDLsyURqcmEd/Epquuwt
KdoixYQTvmEe3qhZMI9c7B1rokSET+aeZUwQ8cyKKmarjLY7fCb3QHxAJ9IyoH3s8wRkNF0AsV75
r9IXWpgaSSHNVKGTJDqU3PXlVLavD5PoTp313CaIDZmkZlw+of+Gf3GQHEaUrsLUrWWASt9v2YKm
cg3UD1BquwNC6/o37eBbwMtCfWHGFbN7SeGEog1hwzad06rf0oSTKKcgDMlpCZMiXTFdBZ1FjdYF
y6MaJ3qLP07U2YAGbJqn2rBe6msuHzke6H58iBK2IXz4hfnC6MEczdP35Q7oTxJIKGN/KpLF1SKp
NucfDMNx2gYmBoggDxnB9i//icVo3dbnYgTZv8TyrrsTRnyw+tc6yl+tldRWAuxi+IkrV011nEU4
euQ19+r0+3bY5vcT+YOyeshoTjUPp049uBuVBAFJlpg5gZtKW5y9OmDxyQ6/g6AT2bxt+be5IPXq
jXcOxrYjzb6q5Q2fQgHR4xKj81Bjmzt8G522AiLWfd09Kor4z9xiXMBW6Md+L6u6EX/Lkj4O+Tzc
3Dj3rETDY/cy+y0fKlsv/sAg+iFLjZrOyxmTK04BDvbucyQGcP2gS9LnhKMxh2WVDvKzKrdis6OT
tyUfObvY8ff2ddPUP2xPcXS9CB2NAWwg0/jH4dIuNVzHK8LBz8KOZix5/88Rfa/n7nC9ofuCA6zs
MwviWUOskkmDspnuxEzwWAwZUTCPlAKPaXB7EfmGzMChpynTvZssPsqTSqhbgeE+8b98RrNMg23k
4R+bv0Qr9YwII5jp4pEL4AbaVN6pBAZZwafeNYom9ktexo6En2we1RPr3KXU9wv2fqUO2v83U8HX
PWlnhVjgsiX8TIWLHiOosBdTswXKi7Yj2XoCB0B7XqXcrKgluto+95easboYecOudyp8wDjiBJs1
WMXt07EgQjuRDu04LkOPY0Z3Fcu9eMCoR/uz5o6uSGcjkisNORcAdRfELYhoGJ9thEZxS5yCfjqT
eRzxx0eDC/HrPyVDuNWezEoOCeXkNHvaCwiqCOGUdnGw3k+B2qGoUXijU9jv++MOzxpTAOesr4g5
vWJxDQ1SSESaXPEmP5kC4BHnOLPef0uJUiBJX8dbPX0KCFYthrGxlWosVsJBYndyvj0OX0Uay4YQ
3tG+gOFykA+0ZJLfVrrFPUARao7d1rViSwA0iREVzQnpeNB7GqTfhAd82cI7ATKa4J5pW8eQf1G7
2vQ3mgm9SzlkOqVRvFEZPqVnDYE466DO8wefqq43YaSxP36UKhnWieNeUym3JXT5U+s06BhYThbh
1STnRdn38FyNhqWy8PXvhsQcFWpfdkn5GrvmZyQIOQ2BAnkLgolFsi/CYLUF9gKKb63dCrRjbyys
Nge7KW8o9sQIMREmhR9tX97XPxJuW8RMzhsdL23Rx3aGU3VDJ+nfgN2ku+LXrZDt8Ukd9KZnfkqK
WbyOwe0DXdyQqIfjHEinrF8KJi9SQGkhRv0Xrnn8U55YpLr4wHV8Tz0xIHtuPNRhwZjBPiENkI/8
Oplb0+LtDrWRoRzs18Jnk1NiMIXAvB0FYyhd+TWVhSm+J15VCoMXlIc26xfUAerOt0xhNVyXgyz6
pX+nj+CK2T4Evsq4yfCAX1fWXLH4pWretSRMXQRYlTDOu9KyUTRYaCvr/CRL8jE/ohd3LyNDnl5a
IuPTNRp4uUtQg8uom4Rvmvx0RRUrgNb3Mhdh+G2pLwJ1+2bnDJczJ51VHZpKLmd9vlwZRs2lDid2
3sYEsIJ5PEwwJ/I87AOThwjqSUBTyLkXLDo3Wtui45vXrh8SCUoXeeEXNNtQqTXhI7l2iEVVxnIv
9uWHcMb45TCTQsQjjfXhurkExgWqMTTBF+33P3vdqo9MGSlaCYrUKxEMCma2x5PMTs6HDCLTDQdP
ugHR4+GUjURHrPAc7ldca2ugB7ILNKtzl7UPOwSXaRidCXV2OdnCbfxvvH//MXOMB8PfI+YeAYj8
zwvNJjtsYhlqhEVY471VoLlXK5y9b9eeSdma1p8xNe2PW7ycXMPGhaduHoJKkBPum19sQ/1VlyBZ
JGN6SBr00FOst2Vo4qamOJX6vkoICh8YOpGDm1TpMUdNWASJ0ToVKW4f7UeCDjeEdv7dtoz+ZboO
j7CvBKuffsac+/hEhQhg/SaThvRUYBLlk5SXGzSeqhsis168msMVbmEQEBlYjGAvCmSwqwSdCLVI
s/0on7UF2ZMU5ybrjIqUXNJEgQQ1/vOYZRGyGFs9XLGum4FgmmD0OiCTfgnMXvQt/5WRDgshEHVn
EEOYEhd0eyFzvsy1HITQ7IxOAneyRRgkfR4J4ADxri2eRMTS9c7glff2UW9dEqzxw2UX7wUcs+lq
5s5PathDF33B+OHTRyVptHak4ugQKUOJmOUYRGT9g3EKTDTp05JJucc4QQ9uUKrYRjPAs5EJoRDi
uHQf0yvbjZV+J1VfRHktByIxWte+l74MNnh6gam8L18ZcTWVlcJW4/DNA5BhP+n5rYqk/Ufyih53
GkYCjniio/ywIx1Qwb2zKJjOqnj3UPl813zOK5C8tAPcSJ6XRTjW53QHdQJlQUyYo+ZecCT0dHN9
KSOZ5HpXXBti6YDpxoTpy50tIZjGTO8lmaNEwxlkTN3rSYftCPYEOKJcEaA7hkSEavma7EarnofX
qvTPX2ceYB2Qf4Glc+UDvyB+pMDFjmSlMWSxzMhPAs4nLPyEZbUpj2GBl1DztoNYLuCX7mESzsbi
4+r/BcbAJ5RPf7VeP5hiboi9ZriM6jx3L5jX1Z8bMr9WAqdF1jXUCdTqlWrU3zRfKG51aw/Nv/VX
EMr5P/OG2Pd6lC4HGrlQxwd9W7UXwyksnpjk+iJNeSqH/6PD2ZWRFPSTf2KgPndE6XgQHJ+c16ay
luE7sHVgP5CuxORtr9m4AOwix6ay92V6tz6fkneBbjOL51z4PXzlOLK/HgiX1L5sAg9yZrn1pw7L
7zBf1feUZYtkII7R+C7kNvsKxEeU900kCBoCeoP1bI6BuhE64izJfpS6nCyldHW9UXkW73QBUpDy
v5h/m8OKWrraiG851L+MAWgLuB3BrufbmY+13/5lBxYEHu1s06nyNV1BRYJz4Mt+TCSiP/72RPPE
E0Mf1QIzFgP6o4DSmz3MYIiBI0+3RrL1y3iYOr049YVLeluAzik0AolhksJ3yQfyXiJP7qRhYGVg
32NNxI/Rwb1kO+wdbSMPxWDphbs/4jjRyVSRyeKDKyMfpEuEJ8e9QFpDkaGdaItyk8YY/i+En0bG
shE9G5QBHJknHvD5wvzc+MM8UJtb4mYox58tvKxJhXhuZD0eIZhLsbmQyi2DhfOc67IpRXrmQHAb
kG7ZPpiJRgjZMhEDiCjnbGfUBxmuIxK3NxkhqhrxFSXHfwAnTl/w02Lw1EiAhxmXk/IWg7xBew5G
8W5+6F8oLvLbCp2k5KESTWOsqtMzqxso5VKQ7Vz3tARRAmQ0txZm9gIukv8jCMmHGIPFPitKJ02g
PB8Tshblw5SfgVDGnEfVShBJ+edmi5L9roSyI2TBfIvAvQxLmPfUpOVtwLMmsCKCKBzpBvnnk61c
fllro8cBuaXmNQQdbwvIGcG6zxvPxMDJM60REWRHvrXCnb5dgBs8fspSUy6qkf0XbKrOcG+ZkJTA
x4SLuqwwBP/fPYHwF3urQL+8rRoQjNJK1NBMnpTvq25ldECsHMKoOoeUHya86NSikd7/t+f2xRno
pu46ACET234mTy6Os8cnbLk2M7GZHq+g59WDfNtUbPkVR4wN9+6sIM4/8CTe4sw7ygXTcfYHAF5l
0i10rmcLx79tBDh/Iy8MoZDLV0FEryoCyQQ6IUPd3bFa/Ax7TmozrhSs9GiZBwaIzYaGGpkgMM53
+kizMMtaH8bU75w9IITX1tx+TZvK4Uhkk1nXo+A6xekAoSvnWbWgtvnIOLncIFLbpw0FRzshj2Od
mv0/7AQZIybORMR6Myzje7Dj+qAaGg90bx6wwQasfEJV5ypT+EMdRRRvsow2xwvI5n4/0JC0cRCs
YeI/s/W4mjbTLSoKHFWuGzwBoSKJIRk2A4sTRicpI9FucHmzdNCnUR5dZhSXc/v+ABwylqbPpyEY
QL9xEyHGcKw88TkAOyJnZhVchUuZpYWG0J23YFPUGEI3pZCfKq2y73sJgELBiYPJJNgaK9uxSFut
wV/6Y9U2sCFewQqBb9ReD3hpAnata6EypYpm3BDfgo9ossMH4Lh+ogt0kquxu3Fjd9UG2WRLXlD2
o7oIFJ/DHAHtwzWSvH5ecM61mUJ5oBEQl+aK8PV4CtXcpPtyyirKTANs5tOo7pf3LkC2QjxcVtxQ
vEUpj7tZeCbnX8yninSEGA/EbNbDHR5Q/khzfp3gYZUzYPVsCH+UYu10AncKhppikI4pgPZDYqnK
o5YyDPckGZR1YLGvLQxusEKueEejCWhQgysl2f+zy3uTXjAbZvPY98K0H4CRFshXBfQnAA6jQ+6w
OhvryhI2Rs8piXw4GUXEAPZ+vq2krXmQTiIbx3qxDju99vW4Sap7zUrpuJs8YJ1HQCt7ypfMglpe
yDdG+NhTyaJfLGeUaH7zsQy5kF8VMhISD9sFN/cIO/Q6deIndmyKzpuX/vdGG14Dv4iiL9XOiBQL
7JC5R2cTqZ66Y+g+QDwQe2Yc2f8rMEllA+iJux5V1+edmL441KZSBO92EIfZlb5W3e8HSWsANN5Q
PLMUTaRdvXqAyw7zgo/hrXPJ+TBPOipTdYCE623auHkHGac8rB6F5nLczh4vbbT7kIOV9zC8Uf/u
UPZLNOWUJO/JCIqnQ6XjWIg5tCnVk5jKQEEsUkaIMhIWw9dLMWuKiHqzbxaE2y3rluwfPQB04hs4
OJSVLVm3v/CCVHjClVzvg9sFdI4lQtWB7b8A7rDOQJERBjXWxl7nGJVhmEdj6WfgpxPsO1S4UYJI
gqm1TBwham1tkB4x3c6342ISOZQCvFf3kSmIwTnslrn18pV/eS7K2usB+EI20pATdniITP6+MNW2
dETskVh3azVyYO4zcHQxGC8BYeSxfdiFExRgClxNTPCL59zNeX+WkeAnDt2b8ro0xdpCKbozyiOD
j7HS74BrpA6U0nZ0cYpPlTPFOgV3bv2lNy0B9gXzveidSdBXW0pB9gE/gWSl7hyo3mnHarw74hDa
GSo+cBUZCfFp+mpHhTWZGXcVjPDG+Rf87AYeShIXXE5Y81nYw4i0NQn4aIyR4xEynwYcaJH19a5A
QI2h8sFoFscun28CnvebNrjcqsRJRygUWQXouhxaS+L78aC+PGM852qBeBXde9MU6HJz2Mu7x+IZ
rI7tb4qma0QdOCv/xfd2SqUC8mD9MAwMMCjclnsVjvkJZHNtczhQ3nYtQMxwXqk29U1jmevcnPPR
IqsUMX3Y09lD2K4Gufa3P9QGzLFlnfOxBu0EnrYRt5TxFHsfg9SNOBrg4BiBddRUr6g5GIvLEFKD
Ei6Fwl56Pz1Q3VZA5A3IB8Xk6k9sJWgLBrpeRMYIQWUCHUGJafdMr6xx58jxkhGzjfL5Lp/fGvHi
3dtR0hijqyC5MBsH938FPikeUUgdVo117nTt/SSS7wp+NrOpDcf+UnHVzgcCkGZ9gVx2nVePw4xT
+xNZ7GRQTfELiQom+GZthQ0QBkSr2LVNuFxLyiyrcdNeTRveaR8Tc2RhXQd6Q8LBl+UlSSAWibpy
mFta/Ki0K0zGo8+3EkKDpN9Op/JVRnUMStvaL1mLjin9zwKptUNCCu6IV1C77EKHs54fbhUZqpeY
P7qjNTTciaLGXdtpVsVcnckxI2R4KhfV1RGes/ZjJfIS7Q20EFou4ZlY/jV8H7She6TqAMF4ClXK
4e8GpAk96P9zCr5MaloyDE7ekpiGoeCk3npaFHFOU4dJK28KRl1vhsb5HshkBNMJ7wY+5HZSvAq7
UkWkqfvjycYzjE8S9k1A5Vx580sqD0Q3Ba+7pkqpFSoPmBRQgfNIwfpcUPjZ6lD+V23u+fULTjPU
tREbycjzYNehdIV6q16PSAUEO3nNYpFxY47GrPEEUE6KSq/C8+A4y1UU1uukj/0LC62M9IeeDw3D
MhtV4khoQQFFVKdlaJYjAW4YtbSUrlSEZE8Wz7oWPWaIbIuAoZUHooZMnW8MPYMwj3tlVOAc9IXC
UuoenLT9OZyQL7Yi/QD12RGUOvdbMOlZUr5N6KykU7PyYQyPj8249ExUkqvxETj1x4hC5lghw5IY
41dHDm61tvtYah+OU9voJaPtglVbWj+CSkoZLrBWXs3d2iG6Xv9ul7USYScFARUSOovg3QQz4tMH
2gIO710p/YXr4vWcG9WGfAkx8Mib6tk3aYEJ9RcM607Hop8cTjPajDE+DgK7loxhF0jYDlaoCnTN
PqHFRQFgcyV4lKi78oztuST+WZuV+y70wbfIIKv5gxapynQ28S8HfP040ZVDKZIHd2wJqkC9oUZd
swqycDs7u1uyQB+6K6PldiOgQG3B5c7BYIkacPBobHA3626DSjr5eQeasUzSnH8glU83pE1ccEix
XrzrIN1CP+NduyNU+ADqbnT2cW6a6sz9n0eQlylIM6xQArY/AoyHU5ebCowXV5V1fGJWalNupxvp
wxoxKvby89QH+2ayE2oZTYUOwM7xJVyBG4earNXT/bwAzowb0VVfMk0mO4snB08CZP5xWuRywpo0
qoX4tUtnJU0QM2Jp/g1GtP5MI8D8NRj2BqxeEeOGlwKmB5sKe7nKwm4/jv97xMcaMpDTivyvX+vf
rqt1gQXaA+bKFXXrJLMkDUZxaYHWfYooaJCIXn47gefWXy4IA9F9UrRrjKmgwwGGHKx5AyuJb+5V
QIIL+A68Q9pXqz+y5x9Uz73roJXTB81mCb2lkHFzOj7IZJ3XODbr15eQndrYJyIND4469lUKXUOz
2cDgkBke8/N9oquW0+lwwT3/btXLj2zLcw5Ek+lSU08tv7wTEbf0U0RvUNYaV8SXSZI6jI0rFMGX
nY7W1pE0pM7J3xezi4Ql5a795nmQ3cFxO3T9cIOoaG3DZx+yagAiGtAX0RMJHzvBBXF/Zt5NtTaI
OoOP4uh6AS4O2wfxI0TP/8PF/SXAvEHyGX7vsWNLxq7/9UMWNjOnvJotFFFNnGBiA8ibBIWnKJZx
pnPbywwox2ZzTeNlbFFWc15+YpwoHabt8/GGODqIt/1T7dQ7G8kgzbq6A5wHd2XonIJJFiLIQk08
XzRxH36Lcx8h2RiHHoK018p4Sdra1wNiLyOqgD55bvS+rRo4N6in6Fb00OLq8xfwp0Bhwq2d2xvr
I0fAln0eCQOflzgj+wpd90hDQlDX6nXafXp5xoN2zX/VcQx8CayUs8JuzyKRgqyntoGfceODxFsS
jOc8zv8lnDd4opUPvNlfegs2KM4ijPdWnJM+dI6Ahy/hNRx3LC7WSM4pWiuNosSZKZv9ncBux5Bq
UERg+5Ll+tcRzZxCgyr9L6Z8k6bdVsVUlwA154LV/6vuHEOvjT8xYB3iNOswWk8osceo4fEopACi
04u4EsIbVy3CfpjqBE3G9XBq3+rraabqEnAIs5HohOIVNio1L4le7NwXbW4G/wL4romV1M54ym3d
IEbsA6jnWb1nPLS/uqGNAAzyT2QLu4dWIb/DHfHnGpMjfc/9HF3pSYKD/vEzKsIhLEgLTO5RQhiX
McNQc/w9gNDCocXhfc3oxHsr5Ssdny7YFlw4RVJ/joPwBzLeMYwTonl373lZ7V7aSs+qYPf0pcem
zIzXSARqlLbvOQqirYUrNiyCU3pT1CcsVyQmoujNHMMLg+OytTJMtutVMiU0Yeo0F1Dt/ArRQ+ST
4XDBEIBryNDIWdFxSCMmjVo2MLb4CGyzgYX4N3Mn5iq6HJC4e0dK4pgGQM46CuYsjJOf8Eb8Kr89
FLcge0YWfxWOZaA8Inl05xZQp6UOyjlpouxjSOVJAwOUNzrDBNyZbbgLmXbDo9uE2f6rVES9FGx3
Z2gUagIHZGJvDBlLTVMn7Sa20vlP/DnFAEBxSXX0594L5cbqs2By0EHejctWPuYMlJ0izb2k8qSq
AnUyn41/BFpLaUo7M8vLK4Boar0VNK9CWjwluHG+J/3440gMLYFKEw0OZuA6JMq9wbTTHntUUwQn
bZ+JuEyGRDfhxhNZ7OyDF2HGUEdmmQoy+Cuo1Lp6uFzoxJM9htWMB5Bfsh2Xj2rbsHuW06Q0zcGo
tsC32T3F+9/R6Ja078fCk+LRY6elV0BmKFQlCfUzXXqqWPa8ay7lyWYQZB54w673S6iNn4v6D+jQ
9Q9vBdTvq7709aissIKJKGpecn9MaB4nZd3sltXYeC3FxbpBq2ho7h0EuVo8Y9zZVbQO6rHJGbZv
9VGlUTzAgWW8ixR3oZNG9GvW2DqQpM4wKGNq+SB3Eo/aM0xnElln7b9BDsGhmDjJx8sEe7y52HpE
ndG6bOUQip4cGyuI9GFHeq794OQCBYMbBQevgrbkSEi7I9SuOiCp2jqH9nhoyGZPN04nA3FQSH+M
5kRoa5G00BKydwNDptiRbU2HqCxgs8oGkRGJerm3A8EuORSObLG4brjSHj5tPgW1kyECD+b2qtYL
UUV1dfjUzIaFlfr3vhXgJLuX66Zn3BgJZLjNHepc+5PXgO+TIkQ8DFlhCAagbRKrmaFTqZRHtbkO
q/PgxceV05LdMtNa6dv+ITxGIIK1DgDT4PXfrHRu3/yZF/+M6BFJw28RndmYyc9gQ6DquGYDRn7d
PJMM7w4FuP99nKsWFfx1+WOQF09Frep1MWbrABGglOXgzTV0rqVMiMan4Mq6BuGJvBSi/6+t57As
S4MN+efPLExlGB1L7mYdj4bB0lSKCDtM+krPPwRL4zK3I7ml/vcmRfgjV61bCGN5KQZ8sGxg1hlt
AiLSaZ7K35Qdp1Y2CZOjrGgtN3jdq8XWXUkxG1APhoFC2AcwnBCZ6g1bHzCpWezm0D8frZTHzDzv
IgiFrXJTz18XxpKkxREwNzap7NHrjt2mbMVVuJDC+L7TDnV15LM9LIECZvpgiZMWfWecioRS/Upk
CWOafRYXaXZfqTTCQW9yxt7dNpltsuV4DsIZvtfBYxOE6BQH4R0NGDETdrv/863pSI7WtcnKCZeW
1adZpEV5qhAFxfdRb1e+Sn7IFvqlatGgRhTSBgj0frwk/e4+QAqMq4W6n1WuqVhp2q+24oknvcgd
t9EyOZkYwjzDthyuoCHYE0adICwlc9CAQYopTBlAejwhAZwz847XirNhNOiURbELdroacAXwebO4
qaP4Y9VBqrbo0+Kqnt45TJy2xnh+5eOwY570rTB2sCXf6DVfWkpM5z8KMu3aj5DCrfp4dp7qvUJ3
9Y2WAHU/f9Lbz1RTjh2ncj2fYym2qWgJkzOninLrBwRpb+xZTJ0ibiVpcA/2/9UHc/tt8sBFA2vn
5ICB/BzDBNlG8uZC5dem0+F+pRlBZr7TuJ5ZZWbPhv9OixfOmLdpPidIO9hs9MqINaYFmYpRlsMw
KZv+1csifhbyJH9As72qbCv6kEBq3chxQHet4tVW69huMJv5CdU0yXKdMErJo6lHPQPzXsw4XNra
Mao8hGhiycSQJl4GSY3JQPaHeIp4tphQU3NfqVZXU0JhdIOlVKDsDaCXG3X01duA9tR3SeE4eTRL
HzFsvGzQ+QwUbtO+vpyRE686SmOAQCFaeEq/aPh2Zxxnf90nA2fb4xNffE+VJKvmnEFJomoWmpWb
RsIBXKBYQTbH98yQiiTPJ3XEEQs2hLNmAGsizoW4v1L/0t9w6uXnTaPNwH8oljq73qiVs4jv+C5f
BL2B6IMgZmptnZVPeEgOCyQI3tnJUXiQOUW7TRDLTxRn8BRnFKgKvnXrqrCUzB1PpEDdaR34pgRA
/jagMWtsvsoh5uXoef6cSP59CeFVcYBnLM/ewTD/AftBmtyIw/fcjiBqmV7sKYno1/jQqReNxpU2
xgDC8FMAbJPT6cJST/hxFj6qrfQSTXm1U3nhWGIw4i83gTJk8Tr5Fn5+edpSvJmSnOixEnG1M03I
QngXnNyDjqafSHpR4SBPaZPEhgR4odpml+ougLfc2HfoKA9trG11Nj3dh5Ai9hWm3NbU8D3ZLVY2
ndIkyBdx1edfRoHf72e1hTAOAZW7IXSD2m8RcZtghMg7/U3VJPmQXOwu72yIb2prRNCMU8akvd7J
z1iUthJ06o5yHVxJvhJoNB6vwG9m7dQCr/Q16A8yTwHRNghGiJKc8DGaCimynUP6NQerOPZNpXBh
vbNi8bF/8z1eSn3/t0LdUHEGzNPTt0ZVuHPDuJF05Szdz/lICTo7iHqxNhUQAQTxoIQT12Ve3KtX
XIHeSeI+7XArHbw7zSuOKqGDmITwb6UNO59U6QJmmb8+OeeCJOgxleU+iCfONAmVU+w32cEKcxjQ
9leq3q9RZxP2TH/r5SbhTe5Pla0tjfIJ9gG7PfogzJ15HYCFiZXrzA/xITzoyGJ/VzrS8EsCx421
rI2fEFxWMt58qp4TBawyHHnWZiqpTg4EdN0B6mYEMhl8qz6cZBkUTV2jLuUjZo03MLvCGJ4EAYgt
x0ScMVGyC69kxxn+4uZ8CfdQ1MRsfCni6ZFmGsbXksilsCfjpo2O6+kCa7XA2dC/PlXCTYIQf8OO
VJTHjaFE9yzEDptYjGYZDMoFdlPqLAFwLf/uF0xfdloYbE65usZUifh+BhYkjhB2vi0PDUBJFoPS
Uwvdmv65F+hGwBjSUmPoacNToB/zAPMQ6Q9zmYHcHEO50u3Jw/vq5EMTc4895t9p9PGWOOzdGNRg
nwA5J5nw+kNUliD6ZBGBYDy23/vHioN8PrfQEk3EVlkSXtYwK5F3ugGY1X4FQ2gWm9GwWHK7hz+M
Dc/6rd/pqeoA+fPre03zmIi5MtQm6h3+BjRsDMNSegaEHenaK7RKAiRzszJhbuSpWBuCM3yzWU45
v3ogqZZC8kbrP7Re5RPxcr1VRxewftoIlgTRmwMlj+5WButUQCPvQfrMtt9/YdueYKwXCD9yNt8l
sS1Jzpnnwg0DYeXrOYaf9zDknqsdZKYniCPr49/pqUMDPU5GkZgsHoRV47XQ8Rlv/yjBVFn7v0xQ
ujCmtS8JF7/4NFm0ObmSS06QRM/zEw/tQzlEu1a1yd//XRgvCGSfH26dkJka1mle3AoRyxzauwW8
tctgenc8zvnrJPoiK1yP+N2MoCGPD2GUO6bSFS10g9W1xy8kD4KURjay23HpzqgdmZfD8+QvPETE
PiiiH1argR4ER0slI4NsoPR6mhiXBbI3ThHdFXNkvHbaa1K6GdVYN4Gf+zP99Xq4J99VPneVWc8T
WL1yiGoHtN4CoAd6ZlJYURm8O8nPXKukrk6tVEknMfxt7oQxnulO75JeAaTDLe3xOywm+F6yxtYd
1y5xCKM8eXnh8aN8D6TH1dhpcGWcXSnmgQ0iTPEGd7KfYtXNwBWDO+4yt15nuzif+xt7iFMhKURd
ryFEzPBS+YmfqRRm7AoGdU6pVNI7QAF6gdADyzIGU1259H4Z3MRuwRvWZSXvCBLghNzv4Z/AY+K5
W76L+e4r7MjVgdV7gXetE2Ed+EEVA+ZOrG4l02BRwx+lj3x7EdvqVcunh/yE+6jNQOC8OQTfVyqb
1/onAWdQPuLScG88/G2FB/VVbJ3jIuB1aojDFcN/AEwoYe6j9NQAMOsk/ldBBHQoCOfsTHOyKncg
6kLyyXC/9wuU9ALouAdF3GAjLDS84Hpxgvkd0wzs6tDXAjeRNPGFPhLkePSozaqhDPwXvIJlb3xQ
zkGZPVn+UBCyitVCdV6P7NiK62vJ2L8QVyS1WVzF9p1VxlgHm3WDc0UDLZ9IucdE8D7IwEh2UgFh
glrYDQKodzUMqIr518U7T5qJe2hVAuls9sPwtQ2OsmHVOSWG0R+Yo5x/YRglJfHOOU3qLiHddmY2
4LMf2oqUGPrNoiB0gWCZ2ZmkFm2JYidQ22nMBJuRQdNruLzfseRg1qLR3wIgH21Dc+Qb+4pGJKSX
cLXvxbO5AMHlpJrEXGqlAG4LTFXTZJm/WsIUGVo7E4j6Vo4K0CALQoD8upq/BpLyX9qirvQgA3gW
PgZAlDI6uv1Kq01BFdMfNyFitAm8MsILmrqV3WMKc0xiC2foDIReyLBNKbwRDgvBrVPIvYkNEMve
WPA5uRN8CvSxi945vlPxfXvsYhGtSCoWwVyEZ+uxKMAMUdCONO6Qm+HrYDPLn86gnd/iN62NEOmf
vEZPVunWkJGQrR1TH+a2dalS6UbUYbukrMwPnwLb3eV/BkPDBdz+2gtbBh88gDLN6kBSJZCpNkJf
URK3bDltKXXNU7LzBgad/zPHp5/0VS7UyPwZ4kMPh239P9W5Dgon03+Hcv0GLce8mksquZpdjyp6
Yg/gztUnYn8COLxNEw5eYBthlO1uGI8hbvzvrLggkrz3UichdDDfdF7jtcTL8jDIDcYQNkaRkBdV
lkL9uRsVBpBgIb7s7Lx7cpSaSVpvGC4hCpbIGzt2WlHXsy6mIMQxJ9qCy+uMxY4/v6YGJHwPhrqA
h82mMMBbBx8x149C2Tqwh4mH8rlpoGOHKhK6XWiSpcbY3cxd9ErgnAniNNMNjJs25GA1qUatWSrj
PiXS62+uWU3veWtQhoxAAYdlm+Oj4OU/C5cqHI7jMz6EwZOGbV32XEoaNC2X3kLpjz2/kMowXcfr
KnhX4D2ZvtmZfOyW2v+nREX0dSpUMEBJHoSqg96Mqi8F4j4mddCIkqybOY+m8gatMx9+qe0byE0h
51+gxwcxUUF6lgtREzlqLcCRK9kR+zWvdoaiio/w2UswRA+ue3k5s4/y/fxoSoNCZbnnHot+JNSl
e3FrlFrswslI2UOrNL3NzKb2vxPjiKOVGL58HxGPbSOhbkLvSVTWsuVdg6myYlgVlvRnc/VFF6pH
YuXbrKDzgjG9D6j9ZpmcFV5odvqCowowiKNJ53hGNApm0Dpfp6zJqbPChQwil2DkYSnxpbDi+E2U
YxZHQ+S6++KSbRiVdV0SmcORHStsV5b1nAAk+06BTJpacvJTRbUmlVxXrMoXYDAuzJAJfJY0ClMn
jO4JzsZE1MCvB4nN6K6lH3MRHyucO1wrXAAEFLy/zBaIWzzIfND+GUVUMlIDYE5hRULFZKi14/5z
8SDjWgiH1dTSX1nxWXqvpHxDpicqONoKrhfvtouPcvpH60EpVchDc11FLOWPwxhaSMHJ6jt4Qijp
wtdnjszYznPo6cMQkKmqSxX3uzI9JM9QNPVncvxTZ6sC7NkfUtQ1vXQz9ebZQl4ZqpHhtpcvBp14
QBpTTiU+lExa/G0b7WqeQ0mcpKIXPlif7NKgVgeGdFsc0wBgpIZ5RDpZWnmMmDBq3cc/4x8tVj2V
CZb6rjDtkrNMCfdFpTTXK0jWqa436Uo3BzA6u5GK5xBJ/H/h5qc0D04qksLjeAo2LL4lobZB6gGK
gMeOtkKxSFl5G8p2HFasq8iVEoxXC+Pvoa8T5NUloTvCJw8mljaGop8w7NkZOAtiEbvBcX08x/dO
P0skA/SpY2I4OhGSvnLl+UnLnrCmtYxYuzByMQCITE2zuuAMcstzcKS0TaVbPj9Bq+Emu6Da7noj
Z0G8k/d8Uiow1cXhTiQ9vg5sVywL8kIsGgYj9tYTjVhvIlSOWlS3D54LSvc/m2fLPIHq2CiLJV3R
FpjdD7BUIc95gwFw0aJRUdHcQDEp146v6ixRLADZpdPwrum2QdMrltQvHpWH9wWCkXrINaNxrZq1
UzwbsUYALlp5E2duD+klJxuD4XI99mPZwiYaAzLBqO+Nxg/k93ZII1g4sbnexL7li5/V7DG4Q2bg
0k0o31ihcTXBtnV5SaUNuobYZaKcoVRNLE0vnzrre1/vWk3HS7rE/ZEWluXyzoZvkus9KVbWLpsd
3gaH9OBPxQVduMjkG6f/bOI2/CRNJeGk4zmvfhi1097IEKYaQnwhTaOHhq3LAWws9L2Z/FsNgjrv
XZQxTY1QftDR2NVLkt+on9WHANNwFebs5kS5CPEdUaadalBQkoir3iIm0WNVuv65xCAjN9keBnxm
QmIZdsRv0sFljV6rP4aQy4FXQXMnIYNS+4MOQ4lZlguSpLBmm/K7LCImqMUJ79aHWTGalkZIgpZc
N+DYmAiTLMBUioj5kZQu9eyt3y7D/X7K0aIkOzLrCnuS3ID9rpEeemaHGP5Dq0AhD5alxd9ZdlXP
FN4bTIlnh+XbC8P/SDd4dD8ftjCcLebaNHTTqVAS/EAM4osOOsitT8QAF2OHJcwgYF5A7yeYv1k3
nI0u6ycbqXI9t0F1qC6/VS/OVlO28+TlHLf3lSggw2uHx1pWKpPpf1WKk0bJ5pOL4qfaTa4VDhAk
FXPH63EfmKePrVIXuCzZqaQw8pKR+LwxOFj9bXQh9T6RPv8xiFi9XrBpaEmwneiBmSfA+WSzuS8P
zVaMoJSRngy5gdWw61SqpzxEXCs92Di4Zjv30QByllfK91WhwD1CzLCewK5enQuj1qVUV7B0TGSC
k+fVrnhCIkHQ9+ceRogT7mCv0PgmmOznCXUszB7TaAcdlobzc10TOV0IWnEeiwGF5mAnpPbJapvq
iUkeJNQwodpKCkXwP1dCisGa+Jqu0uz/ULo/m9tGx2ucq0be4YhjXb54s8yOVgsDTvyXEGnfvzJe
SdTY0DSY8ahpNE0GpZ54PNMh/NxsPuss+WvaUd0o/BDtRliYxw97OBcZPBGC758XOyaUKs6Mg1Mw
OB69s1cvgIb7UL/OuFP9XK6yr9U1nvbHdMW8xfbVfE3+hW/tYLjrxBnlQSY2B7WLSKVCVdWAVbVM
sHaCwK7EBuPuKNmClNZGaLFDLMgOUW1zY/UL911uWWq7Ujzt9KslgSfgCu9dW6Koo25iRlKonBC8
111qu+Oipk5UqGx/BDnH4xVmIieZP1yQOyUh4IyCGfG1gITmTNajzrJ3UhqM7nB+YqhlCtZzR1Ul
yzv+pFKN4ULCratf8RkNZbVnKFHtz498zdrAQVRuGIUPL4trrzE1rli4CVoLxS/MGHfj0D2DQLtU
9Tg3F0chmVIMZ5LTmADnkBX0IJIlzSorFxbk074AgUDzH+ot4OdHA+Cx9UzEEFDvaRVujxZAJpM0
CwXiC/EB7Td99TUnrM6Q3QUE+DuVtMgpHTavFTy2t4XjgXS5Lk6cyHyGhavCCXGacgcZBeUwiV9z
NKSegw3M6z3xgjOHewpn5wqD2aSzVTk6DYNhjh+C8V2TnT13szZuGg9lATkppOa1OyAHIFRREcLw
LU8+rD6RxS2jUrvbw02U2qDhAnRRRJjKVQ3IW7HYVjU+MTKO04uXaAu4aPhXoLm4JA9/PSWqBmd7
62Im6dC5W78vVB1TDlnwNXat7lAPlfTaXMloGmowla0t84gs/7MLvC8b/SWn7mD+lWe69jH+YmiT
yuMinDNg0JAnp31By7UrfCRTCbgPd6zRlKDvMSrLs7NDVNFBgu0PJyKdsZdvmSImWNKKnS3RFt+u
vBDLZhEvr3rGrDZ11wwc/ob4qmfaQYgTKeRNpDKGBBD3fC3ukTaVWP9eD3wcVkb1WvSXCoRYKgvm
0QfPLg9//0RM4T44BZzG5CFSzpJykXCMn8fEg1NfwtYJIP4H+IqoyhgaFMcbYonUN7g7cbiyr5lY
OZrIoo3Ui+N8/MK5Mi7TbYh4PQYj/tAOrBt8Vu+h/RFpvLd/EmkufcRWDfBSSNSOZK1llXv9qgy0
b6EYiTP3Z1/Rz1XonrGcJl3l2VUwx3HS+/6iJLQF5mv4rYXMXabUPBq+gKn0MeRfsxLFu/y83fQ5
TgHA5tqST27sAYSSzlTqHLTk3yRDqiAgBah3D1HlKjqPezSnjOABR2uuoXmGDh39eNzzKXC50Olt
OuLQbToBzZkjDke7l/+dDRCha9zmLEMs6xDCFTYsFYmfPGMkAUCHJV14GFtrntEdTkbulbFQs5h3
2U12kjOFSSYDD/q7rg/7TAObEtTA2SqTKn8+a4F3KYP9YlB/YIwIVfP/6fVbOVL11LsN5+bdGqXK
iD7oIoDALDW+8rXBqcADc2Yr1/4Dp/Wgh+H5A8VeMvy0Kx4lQ1+gF3idihTDqwO5ywrIVq5laazs
0fIPVMF+uSubtQTuqalYTzJY/vCe9mi1bBSzVGxNWDCnTmEIkiAfWxdwu5uB6J1o/PBtO0Ljysw6
fGbBeKv28qrlF1SrtjizAZxB51S76ZPAozkXBAh2MIEXQXia5naDtSFiiBurjtKo7TbfQ8GptCma
CNtt0Q637A9Jv8C7dd/Ph+mW+W684GeJgeJTd+YjTqcxdNSJ7Cr+rynTCYUTlIj9WnG9ZDKwAtC6
n8iM08898IGwSkmHr7DgA4lbWqQ1+W/53dV61kX41ecqnsLhCNiWvnT5Iilbt7lkeb8fPknXPHyM
BkHcVaIlNS3kp4LtFLWHrkWW6/YqSkPK3fMqHFZTA1dYB/LFjri53joAL+6Cs7i6HI91G+uFyORl
XUq0IgRV3b/IRHfXq3+BiJB4El2Jgd75JuVM2kjvWKiicUrqhR4/FFZdI54DDTZLIAV20PAzYQ1z
i6HnyMFgQupGsubDPcynMPDsuowT0v1/7hDLWc8J7n1JSu4l5CxFj5OywrpHhc5S3kx/idt4mSv0
TuqdAb7FSQPp3R2Ch/6kSLw7jibuojTas9EV3VhtxPat0TYhy9fuxdXt3ieRJYYwnJsDlvHyLz+D
EM1vCOLWoElnLeT0CsA+FUkt/TWpKJMQbRz8EDLpRgAQ3pAhA2XI54E7g9VcSHNAaM10yEQ9Ogeq
oyVTlyFBIZl3NLDYTnfaX0GaatUZmxM06ERVZ/rpCuxBt/hruwpEa+VvR/nm/sOUgBZ2brejTKGn
QdM8WEONUWujFbWvBlLnPgOfZoTvvkCGirFaY8SAhQSRvLXyMmytwZdvzlg6R+Sf1TNhxjwC342S
IfJcotpgoqcZfqoV/9rYMCiWNA2/QibPNcWbub6V5paB9Sro5n4Pgac2ETBttVTHWTCDPp0BcV/j
bFdX92H4kR5iU2jeYKI2qFq5Wt4NgoJ0JltonQkAanJ1KZ3HnUrxI/Q45Zh08gxaHJyNVTXiWvmd
PN1wU5ZcoAGNp7n4Rimw/PDZQCkRlZD4sKmbzaCYb/es0D72XmRiha9ZL0Pu4294C08Goob8Sn0J
/u4kzT6eVb0ka1jUs78jhyubeDQ+KFWxDH5cERjOZ5SL8dl9Nl1+Xlr0VfU6k+No3G9qCb3/Y3ci
pqQloBqMFXOrHonwnfQp+o8Y//K45/OFEVBwwz4UBl9ttFoCucG6tHVmuxZeLF8uZ+qRL+XEed1I
RLk3JH4p1OxFMXH0XGTAdThkYxLvnteR2rmVnzuCsJst5xIVDOa1JRJSGBS8qxXyuRJG7iMCNHH0
Tkiqi8cMArGLqbLiSq6oBugk34BduCYq1RHHfCdhTnmexy/kkLByBkllIXEPFWVrS2agaiYFrN2r
onPG71ei4VWfShVA4ELd9UtpkMRwZpZsT1NiAz6cwFwxn1oBn6o7IzkduDTliaOLxSHQ5fc0+4fw
586wNzts17hBXBLhMxIiCM4BhZUWKjK8IKxUFK2d7GKrzdOQ/TUVy/MRNVHnmCLJr35fl9ApKmA7
pCxFP9xz5hopito7kzAJjJGFJ6dqxejLee3z4O9P2wPHWZJ/hC0ZUQMAv2Dx7+LIzsvdeS+j3zGm
dtCkYyt0bTLwCPxXgNU5811cDO5LsA7OC3XmvkYTui9E7SVkDSp6b16QkZHqK+hPVVdFgBoGxRWT
/1LDDUwBLh8Mtff+1hRVo2aMQbascXQCBLqm7D3FubwqY0iPm/iDBvs3pwJ/fd34CZ5OdVCCWZMb
d1Ye5WqgfVQkJN1ksAxUZgf7xTMVe7ySGos6e/C5xVuH+5tlPnBHYR2skDhMoP8gOQi0pYQ+xnpM
s8JJWDhU+1lZ1AsTqrCxy2Hv0HR4ehimrKUx4oK2bxua4PJjFd2rFsxcKC8frnKJsaaKHACQkLop
Mam6rpYDfYc25o9khDt0Nm0jCslwc4kmnYRNy/+wgm0NvLQey4pH+BAgLH46NzTkojhKEWXrXsBr
dE1vGj4WFr41EocrgTP9qfc+VZzTqOTkTrmHHyxRbo5LJ5Qh6gAe0pJWM5k7hibWIR37eBdwVnea
qs0lcza7sZS+/F/m22SBbIpRZGPx/YWX2Wklgd+sG7Q0JZHfbQLVBE8MgaktF4ukZmt0R4eSGn1K
AxqgHHLH8aStWQKnv1M1sKtqznwvMar4kKLRBy4e3O7icjunn9LyuvsarEGPr3EIvWWiyaLw0s2U
V3YFbw2GygHPPz/XIubIrL3K41iVPuiD5p8PZMllKtpNp+WELXFok7ym2UbQiCt/Dk+okAPGQXan
fT35oB2ydPmQ7d/66LiLde5Jo3P7zPLVDZriL4ukqlbkGb/6pXEdWhdGmwN+DfIxmRTB/h7HNReT
zCDPFDsb9pp9cic/8E2BXrWfiWMhSb86HBf42mfG5kcQw/anXiYAwx1YHFfHUMqhijLgqkD9Vt/j
YMOPo3gjsiCfuucNmtVYNqj8TcemazBPK1CWe4Zy374py7fJNhMAivD/MV7YdLEvj2Ri/saGGbsl
IsmZlQ9MvcAxjBVGTCpJPC7TjO0c8oQH70a3lcC3UvvxZJ0PbD9YMxkcn9T0ZHLrDcveupRzEbNx
dMDxKp6jMnU9GifvEnDs2xH+M6h+S1QncFENYMGIFpNEJKec4EQGv69gIMytGcyLitMMbrGrc328
qZdR1+epKfc3UJi9LuJOwAfD1Rbn2hV1twLyv1d+q8SvYd02QGOPkfMGYLyCT4XOCoJCXwBWzkMb
31L3fKdvOKOyJ2MCrDIPXOrj440XqiDF8a3HI30C4Jro6kNY4W9u/JEky3H1N36KlogyxVnFIKuH
zhu6n+EE+5gacmbQOc3Uv9rhKWMHkdWrhiCUHRvlrUxsRpNOEuwxSEZSP9T1egjUIuI7nnVqtbkr
9yCmLjVSw/S3sWnvW/3kwhz9L3qfQiVUg3sJNYtMCtVvnugL9246JnnXH2n3TJ504uAGo2taUWVU
5xelcro32Qk2d6eB+CMLiFmOf7Sz9twRdsVH4fwQXSSRt75v75FyLoux2/Z6VYjLOA+TjZlJwvlY
9YjuXHTttWMsyc7EyNPnZhqKjrqHk3WudU/M+TErrhnHhf4hJn8DOaNzi0iLPYIvE+ZioNooaGf1
GCZnOhkjQkAV+PXbn2WUti62zvbCnKWFZKnkeWUzj9DGnVcXsZYI4pVrNbjjxF+fdAnqW1/YEoi2
D5AmZOX9U2pUuD4+kYaewhIh9888TlPcBlueD79nucWVaZ25+0ivhA4icDlBDbTkNBIbmxm5NSiy
YnOFKWA2bZ5fis/+N7ctBVNJfbAVKz9+/xRuqdRqUpwtnSyHffpUn34ysHVHS2Mx38+ObjxY3pHj
lHdXUaa9ujYwpol3dm5JmEld9oUSPXvnxmRYcDXN3oN3bwPoMuiFGiM1qJ3mbJLUA4MEfPYc1OzA
BmGFkxXQaPTum7rO4zr+XVkstqnW+CekZcXrTbsmKURURAHuYYo5NMVWTRItI4nm34pmDkssAjmS
zurmcC2Pn+bTcDG/j2kBvyYZIrNmWNsdSwl2WLN1jvGflEZ8b3qHLaMJD7t4UX5AJbGNl0E0BOn8
nb0yftOwUc6nim9fLHzAFOe6VxfZ9/vyl3ieQAUv46Pxx3GJgquv1jl56vJ01ZC11pCMHtao+dEv
BGxTFxCfPAAaQjEZLJRiP/So32u05zLu79c66nk/XyyaaiYSmlmBqTOhostZba1sybK8GV8FBwhC
SKelSuGRPskgaw9+HdraOHUyc5lqHHcyy3abrvmrcCnbcz0uVeiwp7e8H4wfuIb9gpomFCupIHVg
PRMMjjPz3f9JO9/MnHZyQuQpTDDyg++NTjNnbrP42m4m/sAdnDrCVXuUcDEDXBhQr4Z+B0iArAkF
j40j5lIJGyZXxiIPpheufv9Lr2pEPjJLwbEpW5gvctE5UAALgoYS2y3E87NcRjl3eODD4e6xaHH/
NBVEEXSr/NhSyDCRG95Wt6vTapoUmNapf5qa0PY50oJ/GOrBgbV78oI+4yE928SVZZN0R2P4UWas
RR30Fmm+PLdpDNUoQDbzXzhZ8PwlzHjeDpFdMC89SscnldfAXiMTPlsmfy0pr5IYFpe60rng/tG6
uR3tTpNdouEfRQuwaSqmR1NGDB9tHAvLHvOuej+0neqpEb2eiQhsgDs8VOWJ2xELZZ904pJuQj8S
Q2A4K7h815szwEqQqIivrGLQ8VAcotRYYdWMse16Gpaw+Yd9fT3ZmMi570nERuy85zbIhVaCG6bt
jXBM4c1dnizAl7EF+Ccfbx7rWGZqFDUKEybOi7tWwfAItpxJkXLPgD0Tx6snk8VPP8wFiBUH8Lfm
yqBA1dJST49z4afyE7VgdbjmF1pQLbmWth2LxnhGbeM+gi4oI0XQbstibSSsgiz8fawltpYfCU5X
//6epn8Ioggi7psDFfsdPVnC6PWU/4sDqzS2JmJBUlNB3s+QkB0GJdMQ0tLtdelK0kYYywPks/I2
638VJN/h6n7tTlxiJ1+pBXXBQ4ksTwY0DxTErn5BsdQdbODOS7kz25/LH5Xg7w/Re/q231GFBPER
zmWJ8AGb+JQeidoVKXjyXJGjNmpobsF8fOnwdM7eY52LzJ/NdTn/op/dYXzTw26Xytlu1X4/bKCm
JhGZKLSbzlE2jP+rib/FSlnknjBzWzpVxLHpaSK7TJcgidkW+1wGtA5s1yIOlfB3MpvM5PGutVsv
L3T4np/EL1iSbAbHt6L8dN5KBmSlKfAIXJq4IFBlig6RH8Mdy8Si2i6YNbXjkXE/QURmez/VibaE
AaHeJbUKaEYc9PHsRLOcXNJGaPSgietCQaY0H1HxRE3gGHr/7ZNyCR9A1RL4O62A4jRgqEMZtGEV
6Atc/ILORHQjwLnbLAzomfc/GVhiZzWBalMriWxPha5NYal0MwNMSG1a1E/8G5LSb8ntpdQfoUmz
/MZpDn04brxNAEg6KJb73bgdCodesHhsO2dvNrXvlQFs2vyUdLSviYfNE8Wu2bEv3LA3Lp4sh9Bx
Dwm8C4NikiG3tltMmSE4zsfyza44N03bnrvlbhFdX5CtBJPj2h+65hp1bb9yYblPCy1g4S3XTF7B
rJcDxyrFw4o7rD3ET3xTEO+OClyhZFaqXC/RLcMJ82pTl7AQNb+u2a3uiYVKggliS/jOcC2tFEuB
atyUVTwXJ2Wk7aJBstwUM4wnc1kgAk/WWI6Drtl6jav8Zwzt/7xexL8FX8236vaVlZPf92KqkWb8
NyLNpFb9JfDhryJaovklChjhX+zS2D7wqDVU1vAavcaxoea2ZGA7+dB2Vdw2uUvjIohy2mIk+GB0
+L6bnAUuJrcQM/ImH9clq53YAq+X6k11kUazzrb8H7gsYJBW6FKgxgew7h28gjvvgXBagF7fUYH/
bn9MISlLtLIxFtu5SINB0hQnH7mflH3wM08TJLgdwgyIMQno0riEE+ObRH9xmN9NeHo1c0AHlhWN
2HkqjQmtGlA1C5vhJbhnfZYVGz2CG/+bxyI7Ltcyu//UfNm+C5okqKF0WdKVEb7Zr7dCskX2USk1
82OE8i5HdmUC1cOGeUrAx5v86LH6oaWk+bhi8cJiqUWRza8BpTEtyutEi6lYEpXwBclmWcUQt+V/
CVj4TsXXH7iUaC2YLnKpZSCb3zvsiVy7jATbCZZZXFWlQX3+qtRIg0yxDuOulJ87Pbnr7XNfkHyH
YGqKz9NG74Mg2ZyGVdqCpyFhK6whyiGohGjbZcbJloA9pyh5MISvTmsT1WaqwMmogoMlnmuRlc/0
wgfk8rcH5txgCWuZ3Wx2AN5xkVAxzU6qf6rxNvD3Qj/XHx+w+m2ITM4DoXr/Vp0QD4NtygROTtTp
wpmFu2xRl4PbJMJ9ZuwNZYMtcmVQ6Id0bysPh+q5kf8rj+qrfejDKmP9AUANbxWh9bB9fFzUo5b5
/H5fuBe/BpFIf0vkZ3ZZ/AZXbhI1Q053uGQbv+XAZ03VM73ivTS252Hfl8yT0O34ZDJUioH1UleK
MOO2x0uWGQFmPNIcVRhIRS5Y1tJohCEho6LoXtKiwonOWr+iMeHsNaAqzLKs7P0psbmUBFjDb7ha
Xe1XzyJxBwrxqHxS5X2y4cqxsWp/j/edx2Fu1Jsr7dJpETcYnbcDbAtVdTcZS49VvJt+2fBiMjA8
hzKf5n90kvuXSrjOwlpma4stZwoXRMSRM+j+Wqsux71DjZ2mOyawQauoAJVdXw++4Y5ncoWunmJJ
Gvfo8PA1MYjslF0091CiB2/Opc7rl9yKELQkjCrRDujxxXdkA6hzYDd8HcN/CNH3t1dQDD7xCfnq
mn7C1M8gjlUtg3AuExHa/ppEguZZ14dM0ZpqTRdkucbKege0s/1CDagOuw55qEU1cld3W54U9GKH
5xv7SYtnGA/W8ziVgxDjj+es4DJa71U6HqH6SgrlpYXpnA1x2Q5M75xY4DM699vexQfkl4f0KSSR
ZcKedA3Ul5/CN5XS6rTklP0/bkkfRFpCJL9DNoZ6g7UG2i9heWCRMa0TaNETtpFQvg7kIHLratOF
eApnsZPZOh1c1dHD5husy9iLnw+ih5lJhUnMChCcZzW9rFOfUGAZQbNiAxTTONnfE2KV9JafZAKE
sdYsBSKF6wi2XCG8wW+azDbs7qByRKt1ROfx7jn9lNrsxavX5jMGhrRpaUvcXugtrJy4/iTDzCib
DH7nkeAsOXYd9YSVUBNB86HmgNGz6Lb53kjBRTV5k0pBcVt3JiAjj/vpO0a4cdKd9HnDz1xrAYsx
/wwKGDOB2hPB2ErQZJvImVnoTUUkNfTl8hxwCE0wdK7ygsu18Nqkd/iMLCAaLLQSEBKmlWOonECN
UudfpIv5bVuiP2hDxo4ms809FKFQzj9Q3LCtUWGGw1uJ/Z5qmcxTtSSPrnkKxo3fq4Qq8Q9N7KcT
2O0pzQuVvfIj1ArWtH0QNvejIHBPim+fS8fXmzvpl1GmxJtTJ+1JB0Xa8J7T8LFGrlAbYIMfHACZ
kTCSvp0IiENTbu4ePKAvbkEDED2qRkTG/BGNIAfYynQ6dBoymObAtit1ZjVhnQCVmK/BO/DAp24n
ZKcAjBEK7uVKHAfW2VS2rsuGIqcnNpC//GgUQ5cZtoMPCUDFiDURVkvniDaKUcuSHBPRJ5ujK3iB
ela4b07S4oWeBTqreH+LaEionFYXVX9/pcZFZh9a5QcOom6nDp1Lf832Y/+vvASoj0O68GRRclO5
M8WMBEnZHa/DASdluGvC5cbCYZ4FbX+kibjn8nwHbxLBQcikVihXAwe2qYMxASTmUQDFUMqKZlOG
/m6Xbey6QzRb72kLgRiDEAM02hPuiiEccrqDw/JYH7ewjc3fNyuInrY4yOoaoDgSqdIuDimSCRvC
KHJrqn6mJbx0/Itlt+SlL5b2qg/WZcFs4fXLG6vnDumga9XkiafyP6BS33pGchuerjelnaobz+4T
p36AQA+w66O6eBsAfPvHdBHhjfMayyfdxwKu8l84O/VmtAHzaj2SoeW3DY9xpMLbb5PWAw7fOfGs
G5eftLus66kmWh6DT7ZP19o77TXQHhaBo+SiAe9D7yTf51eJV1If293R4+26FkA9ulT9czPCfigQ
8LgQk414M84xUpFLdOH7YHAgmhu3fTC0Q610QIJXn1LmRAUE/+FKRY1KzW50Jq0uoFbFyRGF651h
wkhcnKbfIqsPomG5yGWPLTR7oSjsBfj+Hou9tNL7pdOtxj6TDEqq28JyBKX4i1I7ykpfRsB5+kUp
j36GyPno+H4NTOoAe4ilhvNoOW9aOxBiAXXw1/35TNCVWF8l3B2ZBrwMftBnEvKSgzyqmlgy/iFT
CEGx4DsaxV7BJcF3GVrPWPXx1wyhqysNhDan7M4fh2Lq68m5S7VT3FY5+lVakqzZKi5EWLU95nQe
tKlEhT/BAqKjdqoM7TOClgS1Vvj+A3rtoJ6KvjylgUQ4WQ5OYdT8B6ADISXAQ2Hc+H15ZJGUlkwc
6PJ1QFelvA3B7d/xaYPwwevNYc0xcVKejiTZwb9yrh5GMTfpKfAHnhgUvFajXCUZJ9UjAToGMInp
He8Lxorv11v20oU8TYTOupYX8mEG2d2gr346Lhe4D3YAPBxRMX9bOUjM3qpgga5dX9CKio014DQk
6a/KhXmvR/Z916SLuwwEQWrCmOWH9WBp86fN8wKqTjVRiERTwBF1bgvQVGnpwoApoLjXGN8R8Hyw
wGRiGOnvifuzfRQkqWSlVEHGusoa9J0hkMoCc2zLQqlKNpW6cWULT37DhodAW4kP638kkOnvtYFZ
2EggeEi2t7NZvB6Ao0ssGUbYvxsVMsLhLPLy3TceYQ2BwS34p1wnh1BBElzW7lJZQFQpgeCyQzOP
/IDDKWCoEqkbImG2Qf3MswBxcXlqe1CIPrWV3+ruh/ULxxP35bEwMXWA651zTmBKPxr6QyObUwq4
NuEq3y1b1udZb9Yprh9d6RWW4aFKI4b1CsuIEzg2V8ompwCP8AWjp/UYUQuDsvQjHCqN9rf1bFRK
wDoFSwpHiTXj+FsRKs7VIq4qZIKpXCNYBzzfwl0zzp+sXGGQsSJTj5jv1xGa7XGmUVu7+vlKrp3C
lZK4Q8SpKZRnuVu8MH34G3kMu+PkhOWJfWTErJ3pxfHiYWiQXHYH+xDrSEKUDej5sg0YwtMxn0/5
WuJo/vqlwZn0v3k0jkGyX1KUnFj+I3kolOtw2wI/eslXrXW6bcDZb42ef+rPRrd1BpZPB2/5gPVL
Kzih4X6CEPgNXiWhgMleFxAigC86lhCjmlVFbmaIOOmNeUjN3v1Oy77a0e/gLaBCAyRdlxocQQf1
1PBWS/GdWEnNS3knOaR6g2534c0VqdX9b2qaQ0BbExrCRhADAYJnm2xMEWwJsjnB9tBrKGJqsd+S
tz5mnT5ruHAuOWi5nfOp6ulY0u6+4WwNXiHRCDBpkaQP37JnBMnvUpUkjzvua/ycKow1MzoOA90/
84SfqjuT+B8FSKyL7a82WSrsbIjNZYpVxkC1Ki5/ENd0R1FV2ZMQ3DnD3CB++RuaSdWV6StK8HvU
QEue+uXHcpkd461C9+e6azamTZ6TWLz3leDzxeHUX7M1WpSa9J/kiDnPmEas+aVI0k1azW5WA6K0
ocFNm/ZkRVZ0pR9v3l/8NZyRoLKGuGJO0g/TTuIiF357Pe4SmLBKUKj2zXqJOqKisWioDpsBVRUb
Lp4CVdFwIzGzqnVyVER1BLATB02DwQ/McPriqp80cbbA7Whzx9rTQKN/SdvXvVdsHE2GMBlxf6Xt
YqEdDIQu6fYQj0FGBb0NgsiAV2GRTNw9LMFwCCXrG+LujNS9LERf1OqLf51pc7SXESgvkzMR9eD8
0vk3c2mhcm3r+4/dXUC+tF653TMLZPGIVO9I3LA4VG3zx4ZmPhAUyD275ZAGWu/u63B533d9Jt+L
Xri6NucWeNa8ZdZPPr4xRxwKn11MZek/Wu6SYqlrSPEGO1ChAYMMja7LMRqePGcekaVVO7k84+wJ
Z1qsMCzsa2fsyyv84BCBw7XRDev5LXYpxZKCj13neViLcUVYkAoQ4dxaBtZKt7/dq+oX5WwKIhWM
ogJFvTkD14Rijl5MOo4+vQ2hCSgGCk7UGN16z2lPKZUBpDj+acvxJ6jpedm0K0fozRM5zQPur09N
jMDxEoPoroNig3as9JVP8UKVapubrLiEuokk6xLWgi0dugAojsc8eZgeR02BtDpRk92vb0MLPg3P
4/DfUoA15RNh7a0laiNZ97WMQjFbA8nIWNdkQqyUNoGFIsjs0WuuiOiV1KO1HOyGluGG38IBI/4L
1pk1aFwfHjMvXgs7sRNvgQNd7N3Ym0o3cxP365H9Jlw1HjOzfKzlKiuNPGsNTJ1a4XC+8ar/WBCE
nNO4Xx3PRdjW8rN6E/ErVn1CLb8lVmX588gwh50cfQ8ad3xtQpyk2sGsaSrkty37QqGgXRS0nvum
w9QUziXl+a1K+/5w0GLS+ic1m29BFkLZgnnajUiqiaXzLiBj0ki9JR8D2/a0vInFGtjmwd2omsER
04K46/XSBTaTYrI2btinWm/Ey8RMpEQMrSJ/zEvN1Yt7ERbxN5BzIYMqngt5VuXKSlvwr0UAkmDF
PHMzGsgfkWv/r6ANrMiX1KeMOVjSYhnKJj7ET3sLoMRRVeZS6tNIneOH5fP5wWJTE5Q7/e+8Tu7w
QJIn5wWarT7oy1ImnhfjJLlx8gzviCchGfK9PPt7tmySVh4YlnmqcnO7iSCqaJQ9Tfi7lcj/ZbNR
GtT/otXI2l5FJdQcP7tnZaNIJlCD2GEkHK1KhiJvTbdarhVCA71Ea4pzeglw8dHfHzTBJggZY/UX
fKorDt+RPg27wXMBlZK4MTZqK+d3IOUyRNo7GHsl6Qw/RXYJ13NlNGvqE5TzAdjt79+VtBZ2KtIt
EeZMpMiyCxb2EYrBINQrGNmyoZ8y6VSoxKNt/LYNsVOHIgKPtt7N5wqLTHwhxQ5tJskjLyGP985N
LjsjNv5K8U4J9owseUCt728YZ1tEUhX7hJbkh2w3mHayOosrGc3fG0ALHc7RNzuEcTAi7TeHbpGy
3DPk7W+Sgwr0Wi75kzEcI9zjtpQjAktVhkTFLycp34spnjXJnr9ehol3TOn7+ttxQxpY5dihRE59
fmSjJr1x1dYXVdLiTwLceNidPRsQxNGz8Wh9ShUpyfEbcb8ia0r026pcAn6qyt5u3Hk2voAhuFtj
W1iSTWRhLa/T1hdiPaOUU5AJw9DFuL96lBYHzytPiz6r4VkurHgXnKVrHWg51SKwldZ/RKVdMVmm
aB1PDWzgaSR0Mo1xBdeHIeLjshtI01IQlBlp/4uxdBV4bJ6SCcMDwDXG2JMg2JYMkDcpU9xK4xrh
PSevRbK5Ug6SuMfAQupgYtx7SOs7ZXRcq/fAJ8bZjrAOIIGbBu+bzo2mX/Cr2N+xu+oJ3+f1uQPG
+CuYJ0RG7pXirkJ5E8rBPxrvOBxXpJFftvb+f6ksUVRPe71CskrOWnmIc+Cs30KRafi7TkJPiRKJ
9/AAtjA3svQWd3g1uCGLKsbpKrW4aZJh7B2Luqik9PZWN2MrtQpbMmpAAQvo1jOMB14eC8kJNsmW
vCezkAWF+QWNi85qCVdCmy8a/WKmEuNGk6GcYYqcKrVippeCaLUVng62I3fdFX5q3dUKC8D/ik1M
bFVgKrzUc0pJ4+yvEyYD1siJrMG250QwNhZvnMH+UljMYnaEw/f2gY1NYi1S6wuELbItuLpFKcv0
dP7BAmkroZyez7qUqRTXyMIz5N2j1XYnF9+L9MrSCHn5zgQAZo+Vu81rtZL/VRz1murrMso0w1GU
w+Xu4zgE35aLIMINsxw7aAXZmZt5f4ZsRDZnIzzqa6O6xd6rz0BqnCdq0M0xzE4cgYlR9b0XpHXj
QoVX2FYRYYuw9NEBaKybBrbZ6KzHl+BcNMTWoWO5rLdDO9slDpj1T2m+dCcmLL05uQ/cmojKNlCE
QmpCSTUU7u3NeAqhA9gTKWRa/911p0T21XcUpajpe/DkZcZR+glPp7B9MxTuwld5APQYdpd4F8FP
SgFGjWzld5oQ9iS6fTTU7zhsAZb4Pl7xv44t3HRLxLsC8qXJgqSoP2ibf9iRVDge2fqi8uZz9UP+
4SQdH7TueoabIHVB5YGMmu6ZCxHAy8GjH9mCM+3KgamZhMXOGK6Awbb02CoQWf91++cCKAvHIkdl
x9HRWgG5jgQncE4uWpJagDO1rmEZJhIpw9719EiLpi1XASI7CkfOUe3vy0GKC/WRxGm63NubKZLe
9wj684rCpY500YWy+PE2kSF7skEjPELAZAfbe3dSd2w/kFoPFnwis/r/8fKiWPiZTwAqn8Kgs0iq
PCGhkIFe92ycVLVZZrBbe/moiYFMFIPavuFfGEy0moL3ubGaR1OnxDIrHl6cNfkRxw8ePgWtCddt
BM089gLIG5/jnntnWxm3yEEBkcfjCXkK72kaCfclZA3vFktaXUMIx0VDS2SdezEIVYaeRyjB/HlT
RS4simNA55RalqKx0XjwhiB7hRzN2PkURgrGP26tOms7zNQ6JyEos11Yvw9Ub3HxeFfm8TxnKopD
Dgrm6FPNzRjS7NNvy9TKNQgW6Nan9um1Hh8ZgkP+pA4sWag1Z91i6EZsfy21o74jzeyeYYfnpZ/T
bQgF7jSV7SbqtiqA335E1hNkyXa7ljUQa8zORxla7WzTvtcSuNbZc2Uu+J6HmuZr4yaykk1Mwppg
2GjV2hpUMAstcKg7sKKFhjoNDQYRq4AnZsK8N5U0uI1Ohj+bKXBcVnrfMQi4JlIVosA11gduZayw
i+H9L1QIj44ycZjcblWUloNYdLSPepSmumbNhYaUddHfh94jaw8skW+qd0cgUaq3bwqtC3LoGHVI
hP5tnfEj+Xas42ZPhrhTeTviIODEkvy/v4gAZ3oALxOdrpP2kiyqNSKuVpM3WKqv1TrGDl906Ham
KZhld5WQR8bILBYHEwMzlqaDWrByNPqgw44mzJss3Qq0+nLyf4bDiPy/GrCjvB3dwo+xtt/jn1U1
QDt8hSnZuKBX7aYjD9h/g6SMg7MhUUviDYDkma5tpvPeZSXItNxb7ycL+RFxwoX8j/sAZ1Lj9c7F
KMddriMNMQNEjxdXq9ZZq19baux1WD/0eGMAYg02XZYqfW+3EVA36gPluiCmDTpEW2KeinJ1RAvg
Fe2ypvTEXCIqoj1ckr6qGeQkWpKGyiD0NwPvgudeytmxLJfTOITtIpbkFqH/AqokzrCe+WyIb0VJ
/VoT8czyYMiz5/eXxKcIv5YjfL47XB2sxWX1NVjR2s9X6W/MzttjgGUHMF7/ChndRdmPVYCcvmAf
TxcVNGypG0ywWWjFpQiXqF/LTSXyYPAcdpBAP/p0bdxc4nQ1YKRtdkPcOsv0flrN9rHClqLJW0DU
DV3uMvk9MCYzeArgSH+q1SztM3vFgo5S4JcEx9E+pDrFuVqqSAiitoBlHxjLHSK7kF5ILD7WCgKj
jrQmiIi5OetCBy5m7nWqOM4uP5ilrADL71RnqVVQ+USIh3BWV67ZCInhzVM5WAApFAxO2e3yspNN
oVxbBkqVEbbHRA12gAo8QcSJiqiGp3esU84wi610yIgzIG4y/pXzG3Jp/2PaXrzwRTZ5p5Ata/5v
29X+y/g1/gvz7oNft7Nub7Q12N62KEx9v/wqOHXPz/JJJRgTQaXAmClSGoXYut+pgpWl/32Vyz92
L8GBI3b3+U0U5RwQGvcCxth5cQHclObh/3wE0SJu88VuYI+Lc2g/R6qfTTWKjgD0QhKf0Ng4UiYd
/sqXvMH8/NT6gyE+2aYnNJVqYcVyQ1qgwYMR7ovk+sze5nTOlFMK05E4pRk7DnOvCWLd0kf9F1H6
moGLEVr/KZARNmHDZALV3o9QPE5kXPlHiWjs0aiYS4ia8RLmG8wfMzZskRjmGMPd1HMUvOjkCwBO
F95fWscyEmSNLLkyysUOjfXHvVG6Vag8JVzG1gxm9skMZMyt5+XDH+yIYHQ4ddnqr85NcEASH6z5
B3Cymjq5eBbSBqvdNadJDvquod/E7yp8y7C8Y69qJDoFrryV19qQzFTiZxeTR9oMRK8+97+s72VH
e9Qs9kSNtOdiWMSrI1qRBkLcmYL3CI93TjUiPuYrgUp+jbHz7/4Fu4HWO5ctHcV/JDUO508knSU3
ugG+gaZou5VUjvzr9tY2IqU/dC4CLj5hiDzqDjTSMiDsjcSbQFeUAoQ/TWb67BfomeGJDO8X9UlS
kW9dE5ujXpbnrnc/lnYKLJjlTSYHVg7xDMwFeZlne37KS/vUMvXxVBaCCvZPNT2hVQ8ryx7pTe2p
U9X0MqJmWTgLIgo50yPkcJGqAlPr0svY7jlwAfIU+cifgTwGu1cM0hNj2kobtG2PKxASejop+rGZ
bniROQ3tEcsCBzJut/R7WkCbQfX+0yNL74FYBfpCbMYZkJb9ZWyIo/6xBs0mCjaQmhbG18zWkiPA
G7Xdr7B6TKusJAUalSXGuI4PVz64ovut7YH0cAcfoj3VD7oTmgun67T5Qnn1Jj5P68uUEy9AM8OI
jmL6ha88nJ+Svm1idQtq6b5xU38zdZRe2/n4AUO9/eyjr4OjiUiVsHMLOiWgiaMKixfKwiezUrsS
abfWqS3oVdYKFX5S9X4midVjGxinKlgimR/p4T0WZZ9aZT5553Tzp28QJLfTU265Shdh3rS1V8DH
BJWeVbodm8CGz9mtoxnQ8iBUKgyTOO/KEqS+38/n4Wip5kPXML9PeqUMxwf3x2ALSkl/1rW51d/k
w7jFajCt8SH4vLRax5HXAvvKPpz4qztC+NsUaUmjaOAxIDVMOJH1U7j9oLLxcP9WgTEAXFqYhi6s
Spinv8fdBap5ObRGQLcdIJwNVV1B/PbZLYZEAMhDbEHThIHMyg/62XOxDh7vZKf/ZrNOph6/GUKc
c73tbAFEqI5kAbfM2yLT+KefGO0xw3CBws90Fx2VGrufARYPxRlkUVdJ3ryTxuejHQr6qpARpuwO
36zZU/rAiKHzflBCvZZv8Osl8gTwgfv86V70s3ewkoW0wJZssXt3hVGoiuYPKjf+6wBO40wnvxor
LF6NtS7hHR0KSd8wpdPKJjIriPDBSW31mKO4wWMmNceu4KBD3phTx7oeDKDQ1E7jaU21Or9lHirp
UhXWGT0n9IeUsIfXvwpZ1QPNcpucyMOy8TcA9rdTjsWfL8uGcufPiB9+hHSmyUg4gEFz7wf4oExh
L0sgDu9jAdyyIarcxAtDLXiH1fmW/wW7OeawBNyBuHRysQmb7sZhmBCqW+IkswZcg9QkSRG+Zr3x
fL3KRZumPvOC7RuX8auL8dPT6102CchOtJiBejj6SYS5hsTIWD2IPSGlWMeV6tq9WncyJ1zLhC3I
Tq8hYE0LKALs9SrRnLPC0TWuUl0eAF+Q9PhuWim7csHyOFdkKRONjrTpihVw1HaQpBjFL8WMabFA
ro7obNGAFpsvP3ULR4aQadZ3MqwrXqcXO3TDJW4vtyGH53Bou1b7RtCMtmTKOSAevuRnkzFyfL5J
TJeUs1POiW9mG+kShM3zXVmTS7WjZ4cXHKPWnuM/R/GgeCfmW90i5VRu2lR8ne/MbjYHtI4gaVG1
gu8Zx+b3qKjqPYv4gvcyAGaC5vEBOrKoJDFJnomD3IIOjXw1YF7Hd6jUx2Z9jSNxP7nkHfP3cP1K
M7/vSjm+RwOjZUJrJ1UxPmtIVmBqB47KVq/VwraoLhUNhosLj14uKB5h5GQ7+P86IXDc2PIRdTOS
XVV8524v9m09VnCXNuIreCDH3OxzC0OyGdkUj4YH5f6Q4YomuiRud+StzXnx0RaHJhTvjzRNRbe9
AX9gCycY0hL2yMTOqsoJzzeR5aMD9YGD8N4/KD266GD5jOUcxpGsLbZw+hcMpCa+xUcvoE/hOJi1
ZIm4GCFQL13ZCsbuRdTBVCJgDo/ZyT2JgZe/nNbXomLPaTLdY44j7dJDtC8Lzg2zGgmrs9YF5//A
gnhxWSClMF6I10DSpcE7rkn9kRsX8vdA2SSK/AZw3x7lW9EWV4Oz2Atjl3AfEmqEOBvZhxaLsZqA
45hhLM+435zGU6JEkqCSRcLnIklAoLwzYE1RJFiagS25MgZelvt2ZT//KKh++vdZ2xJ4BIAIoLN2
U/18VfD3yD2JEdtGp27WfHdVh8uWD+y90WUYfUxOuy4Zj/EtB3OF7DsrSi2O+MkNDyYvrFGFZw6o
usdy32qzGM53E5ydLKLdDNnFj1/ky/aBJLaHC1TkK9QFgOUGkUgYcduzuIR3B6Fk2mDYQOIiVjgE
/6g3O/n93RYK87E3m8ErdWPHWUqCp5u5CQofQFjwAcTaWAtjyCI3auxKrwnWKibAfMwwUnQLQsZe
E0kxPLkXAc5J7KGbex+zaVFjYE9wS5FZdV2DBh0JOzbTRRpi97bB0bXdf/ikVENYdnnXi4eWfI1r
Jb6ezXunVRZrkifkfdYwHrBhKIUyvtsYEYbzfFq3QoX8+9vnjVZk9W9OHUs5e1X/SH27GxDo34P3
i2CaTC0vkGHOOt5rOt/ipK2ANGVVQbbQf767v5F1BdOS9GoXAro5blDehP2Ru6bcxzbrtCyxPmcB
yer7MfTPZQKX95IfDy+yihGXvLCgVVt48vfyMGwgLFYEVLGSbfnos2VoXg6A3BZ+2d0fr//jV6iY
OzLVv5N+nOrIfN0jzs4twwFQrHaH4ZuzHq0A2KmBe6F4sxTjb/UUlPcixKzRHVODHeqmWloHqMYk
Y70hbU63D6kvSBz/gatIfMnsz3R/NF5rsTX4VJkGtCTapWoUXuPvSZf9ycKR1x9oR3YYySzgjYxJ
BwT3TQAzgYa3EzPlql+/GjqOe1kvoY7AeTSR0jsW0dAZidfuwxkJNwm0ntTpyWU0j4uo5PpK54EL
diAei7XIIP2P7pPiNwqmbwKg8q3Yatm3XCGGIiZQueLyiAz36vcAfYXcH6utm0y8IuZpRItvw1YK
6cY2Xxq4IX4C4H6h1LNG+Gge8kuR3hLn8puxHmSmlQr6qaHfbx0fp6VAuYZsJBwuJMreg2rtYUl8
wSr3rHIcFZG8khlJhJtm8+wNTi4wHa7PeR9UgB/vLEtdg0sNKhG7zuHqYTmdXIGHBbbbwHDNGAJb
Nm9wPmX03vQcDUNCef/qcYCZouYRI5Tq+5OaZyLGfzA/COXMgl92XlxgcRrOODr329UVW7qOXYee
ehWTGtxvgxfE5dGUDz77KLF+o69aKdWUYT37+ROZmcDUp/ZwfljjquY0VVPGNmC3ELQ8W1xEXDAk
pm38oxdSnoLVQ7etjon7GKgG54vUvIkTEx2dF6C/01qQ/bg+wL9k15XFmcMSFzJNR5qnnm2SRadF
K3kr6FZVWDBzyPX+0km7mUFbdfzySnyltIo4NXEUip6aygUCrtYngXNJEKtshxUd+90/DL7I84IK
1H+4FTSkRAqUWOIX5nxMtLN2clZbvTEvPQO24keWIo2Y2JlGJgo11uHGS1Eq0QmamM50Ia5tTNVv
dNraj4eFtDYL8fz6cSYJZPNpu1gTGmtofHmb6WdTutr/zm7jLmkVZWqwPLI8Fai0WHDY4BfbzUEw
c2+2dt/5mF53WtapgW041bbfBtIVtbQMYIa7wEArIT+9oMiseRug0c/tiZwjILNjCdERn1Nux9u+
ecOLLNuhgneG22liubzdlUU2LoO12C3GFOwnHrMMvBt+lepcN7c+dVv7CIT+2y2wclw2YpVTFhwf
tcIjbFWBBbiO0JYQAlyxgwH0RlWUvkaol6NSrG2+0DHR0MA88w87AvXxR2IzXBwUlXeTOeRRwBj/
JzWGAmtoHr1qGTD+JqE8fIYwc6+WLGgPqrgdmXNvAa3EviK0rlUI15AaXgcrheNDO2qJAIo1bcJ+
5C0NleodIi4iBxd7eRSencK1AhfY/t1TM9MTKb16UnZTRFS70I+UcITqIlnuM08OmDFVWR2kfX1+
po5HlH2FazZCPHBgmT644B1jkjVrd8K2k+WwKVLB+XrOtB6vcSfO9geVoWb5ObZLyLNXxmunuRqL
UxEMp7Snd/pW5COjczy4vrbc+M8xXvE1ZjCuQbaLVLIT1fV5d83fjcO8fgpIR7KSinkLQduUPJ/8
KsySZQifvHeQegvaaxBZKwZOX068xw9fzIe4Kn2rwNyAMmjrNnnb1jtzZwU1z67lZanUaRAEivy8
6BLYKgSU9bst6LW91w/DHQJOI6AgqhtM5sG9fDqPJw08qFa60OAKL23Bua63ITNH32JmvbggRsJ6
3ydnLuN/gh8lOK76uD7uL+GiZhNu25FdXc3dAcQcKER4Rkp1T12wj0wOQq8IgFoqrVKJ65zWiBLF
Yp76Hum+8j+7EsbZRpAmuAk3tT/NYivfKkK+M1bLRrbmOVWORyCCldbh8cnnwvm2DA4jOPuGbSzL
r7Hvt1qnwSOEm+dOHgNVy6dmzL+RO3RqbG119kfk4caccdfmn4FWyXCRwXgzKWKNBR5gB08HFMwS
eNlko+uMrz/E0nHziA0wOFb6qVrnqAx2aB3PcaoF5+tF8gut2dUURpp2/mkWiScF1hPX9Dhbi4Wq
/9+mr3ESYuMggaXvXwRGz0V2ZjZGbped14V+AZrqtwlyCyGzyHAacjh+7EfSl5Bz/otAY1sPu0Dr
5NuHnlaNmfeQCiSXG/8D6cCBfh/HUjPGzqTqWROnMBk7IsZBpkGDU31KXEIrnQEJiPui4ltz8Z43
LbifGusx6wDgxCUi3YbutorNZoTAYAUcU7lqU6p7o46bMLD5UtTeDvQvgrq/wEfAmfl4ybUq+dlF
909sirmu+5GL+1/eDOEEJx3l4cFpYhiUnvLg0Wq3iDGSMIMT3m18g9WzHJxDPpsVuef1ZpP+WP52
x7WJ/+gSS+dc7KIpsMOwFRc5M5tIDytucGQDrYdaFw2RANo/Y+DT5c+THhBFPnGMsx5QgkuOEqI+
oebXP8qdp7A5fsR8fzv4n1xkakqYBH2XbeluGFOCGZQU1tfyOclGJckXLjMWGEUTg8ysiYeOUmju
msvutERC7IWvazkbe4/9fbK+mfFSc9yoQQPs5cZ+6+lf7WWYz7++ygeh3Dyk0Fj6eWuaA4XuK+mT
3q5O43PkckT18s5zHTLBHOP4ZFjCIkT/1J7V7LUsmgmoC5F7zC/riDZkEZEEMw9NzoTmprtX3QPg
F8xwlZBT1ZurgRpfqUiQlXp/Sy7izcJV9rW3u4hlTwQRcZdyz7dVg5hTL/fnREAP9YHIKU4BMdj1
6tFLX2PNmy0aF8emzmt+J8ZuX+DYAyRpN7LfhRd9WZdxuG0yuoG9oqw8EHAOf6vZUb5HFnqHbdRl
gr1aJKQRm76NaKeJVxvJfyrkRrGgXPzTuCL1Zv6+zIHeWHzhQPRWRhMVzwvzUJBnMOnPMJMmPo9C
vFjYAHDi+v3R3Y7gRxkpuxstXub1M641Cc9GYlRbMHio9MA8FyJBU4CfNPD3dpTtkyddLy2fpTY4
sDLLgXGyNB4OpDpK1UY2OlzQ334+NHbx7YjwOGwaaNBEP2ftdJjvkynVnO0vLyg2CbXPwSwq+XRK
r0J78hQ/nyZjAOVakZVoUacFCH68nAeEvPjv2pW/ssa+RnA2q1TX4wHWJjS4fz/qbIL0vZt+RLn5
xcU7kPbYXflD+iRltgVKYlM5uqWKEf+7m5qXrI1KMxwOHxGVsKvmhhI32gpZ9v9zyCyAOESt/oz5
X//za9qm0YaXK4f8SiU5fnoH3nuw3MEQ6xAdnEoiroImAUJ6FQkgVBu4IoVO44m4F12SBpJWOw87
yqgY2iF9fCru7tL/IIEnlSbJOEOoc5EzUAQAb0y1M4HLC44Is1X73SDH2s8y0bK6gR8A4ewCMeAQ
hy7rWdHkw/nzrBLr89ZA1Fd+UU4LUoIlpUnSed11sk0e196yCo17PPNwAjhJ5YXALeCaEOfGb52W
Zlp5ViuQOL3hxHQ7XqZRx7a6Gg5lBMF5XNb/Awj6075XnPMVWIPKgsE+nFQqzdnYwneCBz6Gi3og
dRatriJYPd9EfnS4ymP3RS3KjKvRf9aelbB+q/Ra3UpdlgFLKAgsjPa5EY8bgRNvhdB4aSdzkwU/
mhnOxUJyUrwCoICH9U9kU3mrXvuPcTTOndbzMoBGoOw56soMF9ClXCcnDZ6OVDKgpaaGO3nK/Zi5
LNJU3MVIM4hhMwT+wMJQCAqUV3MpbTCKp3dveitWNYD10zU7xWlkdyR1c09xK/G2Jo3KZM/r2wGH
Lpko/SvKWw0iB7rHJ6u3TKkStBoUCFZLvZPFgtuwEr5fTIdi7a5j4JONVHSUxCCb9S4KoLkQ6Hiw
fJ+3uFjUQIlinmU9q0OOx2lE/Zy8yc+ItPNyGqquqiw6ioLFB6DI/ul+Au1bKur0nOw9EPwQQMwi
zvfcjwFnMVDVRcXr4YcElcAgKNvTSa/dAcFCqZhBVfR3CWoXNQC0fxO16J9MtVvnb7ozOEUmYf8T
yWaAh960sN9MNauOb6AW+J8d2d8GPgAJN1s20RXijlJZFj0FXCWHbLagBxSDU8e2wga1craUzPg5
PCmQ0piGVcdIGzCdcLy6WVBfRw+cPd86zAySvnW1Gz5BKrtJoMkDfLdbJE9iTmV7k77NyJwOa76+
LDaHWD2eA4/TxVkwdFKDGrtid2CiJUlOpeJZbZ0Mm0cYXUTSWqwyVo3bIweofrgXoN73oEGt6OrT
3TNTKAf2cDKTraM9BGRDaQ/L1SSnRq5QMwuQSkpPbjltgNY9QJrUkAoBE1PaaJCZWClB3Au8oTP6
iF9uBaJlUYheb6SEwCCxWKA84U3iPzK7/mm0I/bLW1xCtO4W6jmfEywcNHlDJEzOSKL0IXsAtblv
iwB7G9ZvEx5duP+/60RMT1QdRhbVoAYXLpwqxf98gU0j6+saSlC92OILz45MoHhKDm+GPNFMTsXc
go1kKGajaR2KxSPJBV5nR9EUqsNEq26hpu95rafpR1cHGiz29OEuhZ2cwFOtTY6aVb5ass86ZH3R
Mmko/Z761gci7/qeCVQh2YJISzGERILN1lmgVHFfXnvOuhZmM+iDV9FvfdVYkvekKg3BT3TfaR/s
EmExLxzeV3OcnPxUqeAHQw8Bfzi/3NtPGqPzTipCT9gQ1hB9sB2lDt8+Arbql0GL1e/ixg4T6Fmq
CTGEPW3Md/7EpcGceYetJ903GO/tL9Cn8U+HjqxRHM8E7z4oLPAyybtZmKbQUT1yQ/GYXl8J2ZNw
Lc2rDGxwQOvjdzH0U7G/xP2wBu1FqJxsTGAAtzWgs+5KJaCRumEWnUz36EDs0ZAiA+IbBf9AAZS8
mhl16lYtP6wJ9F4SW1ydlDv9SeGRioV50uNVCQehwIiCqXBo9kqkpoSosCCOkvxXXUclteqW3w64
R3VTsBzP2kHRwoM4xt35AgAoYcIpzZesb7eVjIOQ1iqsRsQHeK8oUUVmIwvPZxCwGjQr57Gy489d
sNj9WRCGosAcUfG2/6kzYgdZee8UOR5225emUDcJBY5aa/UEoIUs6hd3a7bQ7HS/FJVRb3c5xgBb
gXX/mvUqJjCbe9rqbZ27SRqzzYq7EKvNgjxH/q9geFX3Oj/g/J669wAQlsIPKTjv7fBhHHLB29yQ
vD85/M+jR6ZSfkmINGleypwxZmJBBLi8b5J7r3K9383wl3Gfx8DMPO8ZFMRrWXDGMi48v+gO9PTp
9y+1rlo9Sx+5o3BAsTbfL3W4Vwp26aH186GhiFpe8UiUmWbbdi/WAaAGfnYqlyXbjKKEQTOy0F9x
7OJHLweVZ+Ib6ehfVGCvcj1n1zHHh6g8wjzkDyPtsaiS3WMpdgiCj0s264sx0XoTa1IAH0tBAH+X
2SPLZ64EA52ZgwIGdM2CfI86zMiVqzWCDPHgmqGVJaunVfCun7v4zkjK0Ei1qEDM98xXBnrrD9cH
vC5Vabyca/aDTkPkhViY19Lg7gqS6KD4bQCDHSxTHHcUZ/Awb0E7X7CBp4fMv8eJGxsw0P1xdT0t
C6VwnRVNgPgi82QEvqPdvKIjEKZo9l/B2at/OV9GdSFodcCrZiN4ARVRIgBmrMUBSA45TAa3yGCc
g9Dbga6C5gTJdCFzj6W2pgZSa0mhDYHvwJ7FOSL+FzMkYcq+LNXanO9raEBq9PWTZiEUCMVytFoG
b1utt0UZEH2SxJ1qL+/8sDoK86DAOu99cIsJMprYPi8ITR8a2MKdTxZsQCFg3QMSwr1Rn7VVN3yB
j/UjuqqklHPg8QSABz5dU/UOU79fi5gUFXSuOXQ+/VlYPtQoroe5dTLVTDiIdxAumfG4jFD4aNSn
a5jNJ66dajLr8SM2EDbUPldK8xWLdiKJOdfnxMKPiyHXJXAkZSZp/3WPt0XCSFP4X6Ssb6SCkHb3
lu6ebiRViUQCV0zmzx+zS7avgL5R+cjrgmIbV6wU5NZZgYf4QkV/6kAnVcd1agYID/A811yZscLR
kAQ5kR71TChvnbxRL7mCo8grY9R3ZpvXpxEpZX0n59haejbrvvEhMvwE/sEOGXHEmFIodqZjaO/t
++FZTJCXvqdbLZQxcEA6ULmtwJbo0IZqDq4qFzM2C9UyOaSMi3SO9c5SIM8iyzkwjISiPp9zgKcc
xgIryJNzZZhP0cLHmJdrgQiLmefcSQaaOqhxMFhUmfJJa1gM/2aGMJC7j+zQgcLar119MWDkohso
9kEq51ljNxbRqrHSLrg1KtyXBZVgzG6zX197rv1LTPEM9FWEaV+OFzgcF6c9myj6r6Tr5ePCORl2
F2bvPSgp783cGOHt0hlHc11D6IRY25wivnDfBK+s1RVK6LUL1QmZHPRjUBuH5Jz5t0yCFdWlntMI
7ucQoU4SKPE9md1dHznouYNQFS4Z6TqXD+qSfh7w8FxpljsvnDKdTFU9CxEbIFOrDuw5VslZpylT
jP1tYOHOhgzTJ+2zvoB4BLoQcP/x8LQEEq/Wv3toeOVx3w7weLMNW8hA9Ge1fkg6HJqQ82APt9XB
p/NCXz5xWmPSm5VzN90uKwP5lImvq8i1VDFcdoLlI4v83vDue8oJq7I2u9+uQnnnBkiIJJ0Dh49f
nBnAf5JsApay/uYIKd2ck7W/tKjxmYM9DFFgz1iSV60TisP6mqpSl4XQ+29R04n/J+vHd0dA17xA
B0qtFge8ZyTnVMQ9KFtrqZXgpGdsfF0mym7HfrzfVSgRGrC/AuO+5bmEUvgOoFj0AWQq6WM+W+pF
6bGFffXMN/BvKNWjy60t3/uT4Ge5/kWzac4wrDyRbbTDHG4MigOyU6Zz5pp5Q8W8iJxY9DtHxzxz
OLKmkfKFLFE4GhbZ4a72oEFrHrBbU1eSFr2O/c+hoGfS0Y1NdfZMM3mU7ZncP00Cj/UWIs0GIlN+
/FUaZ0RZcRPCmiQRgRJj3l4B8sYj/A03ZJ8FJw9wqJ9VleMedBhdocR/RbaFjHbhrPcjFrkKUkKP
5uTHNQlu6h+zLsnfXQx6n8M6NDSrJwYrVM7+OsGPY+N6aXcD6p4WplWmLP0jUKZKJyNMvELwDRxE
J/vE8cppB10Q8KG+jeIpOquKGmaNSUw2MIJnA+pzt/mWCWKRhlrOszhL4ZaYRs8BKCDd0rUJ+45N
+4rj4Rbcnk27g30FmJDJyVmiX/sbGVQWGxo2PI9DbxeKYNIZRd/Ulc4JGzNpUEegnR4nHtzgJWIW
XAOm8wwZgYRR4WtEU2GKAs/GglcdAUh1AFh5bdI0+gHfLE68uwcMp7h9Uie1YFBo9X1+m+0MUN1M
zGWMBn1e0gMcTNS5T6xbA9e5XtrR3EV0O00mBGhPrskC1M3WSq9MXQdsRMBLwPwHDysoORDfeWle
iskUoHBbbNmsP/7lQNvncfw879ONCvCN71ebM9cxWcgR63UdA/IGOca44PRSa8dlYBrJ4uhir76y
KOOfkFFE/fLAS1ZRgwGc3lBEuaCu5cbfb6aLWqKCnVy/x3bvtx3EQx0AmBBeJzvf91H+h4BCxssU
B19JpWM/yV8mDD8GjYP3vXU2TudqCje2JtLXQmFCzpUBlJzR9v3I/zlBlsuJ8oQnS/c17rG3GMG7
43jcOzGvR/+sZ6riJtMp+Oe5LRpEwsw5EYfwcMKMiIK0hGA/IANIZHJUltzVQPyUJxahOED5Gqsu
+o8pRDazm5K4Q8y3TLBtgDQXn/zK1pIzwaNp7pQeFHwpAmBV4Wmih7lF8QIel0wguJddZje60gb2
+IOX1RJlqhoERFbyrsmeQe7aRq2OhdO4fyGXLHaxGFRy9mIp8b5o589G/kUedRVCd3NkOzPnelPZ
45yjkVjK8VaHCsCOJ3KlFktet6mB/FK3GCRDNuCjljxlM17pyR2mo6t454UcBCDn/reyzSgvOXvs
ZTR2DgadIXMGswAqVMlkh+n6FH6nJI2G5O858+Xr7q899kiOZIk3QmWkdVkyzY6/5eH2s/KZ20/y
xeRzCgmIkNr6cYFuzP/WyI2uids7EmwYa2MjzZpnKpl/7HENpFEBkrHAdqteBPdWAPbi3j9QHI42
sbE+4L+OJOGxVP84dNno/3edU1Kq5dQNRxQnXWktSwc7ASg7nUZzmqfA4mhEhp12rDmrlzLrXNIm
GhaF8QXu9zBd90pDwrpM5UM1W3Zbt9OZSBJ9fE1354v2Hm4a/+YGLPR1UznHBAOTGBB2+fs9pjbh
P9+vhf4stzeXEnUDF6tdJN1lEC1wAAR+ah1T0ukAvlayQQz45IEKVPDjptfHGYYRuLxvGSQJrWm1
NF7yhcQ+0jAiQclLh2lAqcykX/9SbPwBT7Hj29YS5kuUb0dpR6rTq6mWC7sxi4/i24zAYcseu9Yp
f6wJsQOmqP7I3AYuRrPN6AS5NWS46oRNx0PWDkVluP6SkNJdk7p/5gPc1fP4eBNZLPvQFAopcONC
jZBYoqJ8cGLbdED6GfnM8k5gCLCoq1koDeA0phcSYU0rM8QIfBV5k0akvyB49yo43sZIMzka7CQs
bFrLBDqoy7akwAV2FZrRzTZ4+Kb9+MynO0nq+zpOhICyNHyRHphdzGFPOWDXc7zb6zw4StzEaPfa
OgVilgkud7QzexQg7Uhl1ZMeO5KxqtOrgdTVtDOKCkbW8I32m0rLQ1AsanO3qDMUp5JS2G6rmo9N
w7xEO7QhRc4rF7zfkXeHy0p5hAbnOb9XkIxVe+XDKDboh7Ngbew2oOLWhWJjx5sOKbMbhW/VHrjn
joTPtpMt7IODrsOBmz/5ygIWimoLcwUEz4rxS3RPZcrxkCqS0d8GYIW5ZVlYiI5LDOvFTs3njLV0
CK8ijNVPbq61g6Y1PkTBQdnQUurBgF92T3pXjfpj3QQJ/qxowl+D5hIUyzFqxCvh1anYPi/zD6cH
mjhcxZ5PmSEDMCJWMyXBk8G9R/cug8DaNyyPrb/joEBQl2Z3B8Bi9yKt6yFffIIoS2wfXdZJ2afE
urleuawl5oHWpoWNQQMwHxNdKmT7CWC5LPbV29OM615JWSGrGX6rwpOcxeXldpiywdcaILSkXgj8
f6JEOlBRz3lkUwA5cD6W1uLuqdQHsuEEoEI8SVc39RyD5KuF9b4GLBSlwPb0Cp6iaFru05wpv2MB
0ejsChUqf1eFxKbMusuisvHLELSrL4GpzvdIQ3fti0bmhVcdaAs4H2Amzr2m5GBBD0M1Pam8GeIh
AMyr4wlgppQVbR2zbAqasLRjJTt9YAnpwZ/hinHNuwIUeYNWIT4TR1MbM+a8foBki481b7kTWCGL
gFW3YYAgtSBOOJ78pI9ZmQOmIXGeLhwmUnrU5pgGAi/mmJDaZKjjIHWdyBoS5sZcwofdMhXww2Nt
4cAjZqDVf4L88lCBuUcJkACzM88Q5w9HDDcprSdgBnY/3mMl/tzMnp6h1/Ey4sr/VDwy9fsPq2Db
yCX7ndlAXslUU43GZKyY7dFxOZrzpHU9ZyUNet+9N0B+U8plyxGF+ExixdyZJKctViuxI5DJJbVc
KAL7NhVhpC8PFc9H5gIJu0BiSejAJ80ezW3aiSe1hmgDBsvgCSOeS8nPwnEWF2l6OkGt+ktxTtw/
pgjF55bTQbrnnyux8hoKNfEWDci/AnyMA1t1Dndqbj+Ic9a8Ci0l8ZR0pR2MMReNT6WhEX+GcOh3
lfmGwW+Vfzb/6J9L9hr5/w/Xg0l38uFlcrTBWLXKXQwb54F4qtmYumQhUBw0MysE2dDNereTM+2l
Aklp8ywKLj0dPCFxpj4EtKRpxZVNpKlJSaFLxGJuRTrFU5LS4gXDsUMLHiDh30gzHcgOt9OESW9C
BvLUx72NMMiyEDxKkByQ8Xk4CCutAoyHz4DPqCvMd279BVu2Lhnz3UOTZXHFfHlhb3f3MUl47+r/
X7ubC2m7bpCXWGHQujYVOZeVFSxv58YCxiHbIfP2K7pr5cYUhpM6ZOqGY9mQh2lSJcDVsPBFBp7V
4hUTYReWqCrAjLU2D0JNM4bMm/refnwoo45JKSQjlbjrKZjbRl2+GZ64bVVddIh8VtkeDx33piTt
7z3awqdMlx+dljAh0C54I4yVy+JN1trs3Uk5VejnI9eRxcePajJGaaMygUzwEbXrQ213Zi943KFf
TG2tc9Xu+q886q4PA6h4/JwNkwJW8jxxUIPzcNJv246bH43MtR/0qFE7P7TW8taNYbbmCiRKmHtE
B9UNN3/+PZmUfsD+zDeo6FCYk3n2nuJXoktR5f3C79yLzDXuUtmIwShSF+J1t/Eir+HJHuuYtj/l
2r6TY+5DQ2Y0kko2oY2Esu1eXUkqPFuwcWMZtPn/0nrm1MCH9gDDvLyGVMNFInVvZ252YFy1kHrt
kukcFER30wphMBpe5kMy8KpHEK2AKJS1SqGXQGV1bK8P4iTZ4wDUldmhPMDW6/5XM3gPjEX9RSLU
XG3W+8Zh7u3Xafatm0mgvpv+51Q0jjwRAekPlXhdq4gvbKxeOo7kCUNYigmwjTq21dC8VlosGZQ3
daLlrq1m8JpxfkgIWRfNPtlFRIUP8TRf6bJ6qYvibAplhSpcs2ycBaQsqS2Jf4PSy9fewt9H7zst
ElSBG7aMq+XkE1RMiRUrsdhBC6+jQC/Q3ESQU27j+FIjYQRZ0TeYHHxxXOJGKFuaegDYz++/PLAF
dvBguCmLdaDzb90nHAUJmBTfU6qo0uQraOGZ0KwsCajoRvM3v2ZRy8ttJ56adJ3h45VgW7sbmJKS
oVzQVPMm0Di7a6aRTJ1KVV5HIw3hSQROQYhiIYQ8intxZJRp+gCm+pqWbtQSvkPofJaBayNiyioV
3soTsBHHema9Hqrih+ppqByNFHGYAfKf8n1pxacCOBBD+xGz5QGz30qFybaHY6eI82aycDDzyaAv
+hVSUbhe79pIA4OLRimJnscslWWitBA7a9qNaOy6N2I8h9+hNrv0e1rH2Db9SO+1ByL/Jy7am05w
gjlMOGo3Py6JWS/pLLzWDFGPFW3M49GtX0xwezD4W/a+Fy6rWMAlrnsyCYfdeOgw5RvK5YhE3d1o
uhNHlgtpTFAmLugtjJQZ4eDkX7UapzER4n7o3Ih5IAl63t6cSkQB/4OYtLWrSzH9SQL52bvEEv2+
SZCFZgnE4y3ViGUdajAxvOxGS8tabJ5oSbRSMdYz2frCUkqXCy2hdHfaagN+OpZgYYZU39nVXdKv
fToc/tZZ8WH3YC/ddGYV+uHPR5Gctu+ej0uK9TIHlqSnxvyQjExthtN4bH1C0HsFWRR+Fionkq2R
FK9EvhI83UeSa0Jw/Ho98kqKQqUjlljbZHO+Mb2HnT4uGRjQSnd3/piLsqGCbTLm4dtzKMFEltTI
KB94aFsc7hnIGlwT9IfNQU1AsrygMEEgwkj6xFFyH4TpFGq+38GogOYDFwd7jrzApmYfxonrktTU
AftaJ13Eq1h0R8enIboZKoYzspE3LSE+cMmDqvnOZ1AQluazduyJJOl92VddGVZIqqJaPxe49PWi
vKmNx04t6qQiczf4ggvBXRRv+5dopfpHtRrxRZatM+xBWby2H4blLOh+AxAblFtdy/vk2St95pEA
iVzUfeCRM8rbQJ+GNTAL53BfxdUpNe8sK7sm25hZ2ap5gX2FqAtHHBSczdMi8rV3w9RWNGRe/I2K
B0bZ92j/MTRkCCtP32ADx4mcNPLfX/F+u+LzzU2nYouLrdG9EflayJ4qsmhFUzPUMV7SAyUfmPus
MXw/ijiXZI9uMMaAt8b8PmNSd8H+nNjmAx2lV42KyCN9ZM1XexWvVCVSwa6biKMLwQ/9xG+gmJ9u
Bsd32oaOiMLxJ4LXVYCvYebI2H8waYjISLYv4RH4Xrb0Gs/HGudi8GC6bqyyyB4/xmYLLOMnvMKD
e/P5Jj7jM95ZHEzOafCSnaFrr0cDkh13+a0v4yVmsr9Ick9i6V9chSCE4dldnHuF0l82kUlCfEpq
5gOmvXFwxCW6Khx81nChjMr2HX6r4A9CKZ5cUBHxEoOjXoSh6oarqkGs/N3kPznCuxsuAyRProEF
khfDJxnncI01D7NlDk/dbF9YwjczSqizYp2ZZaubbInLO2UDTV77jKVUfUk2jJfc0rDmR6HK8nXb
d+BuHnCFXlpJ0VlvxC5CwAafcGLS5hpRegutz5g6P3U7AzsS2BLXZDn66Lz6V5VSQ9ghdLAOPszh
OXwSkGG5PIb8KDPXcHyIQWvtwumVIuZ47gwlRDn/bzi1sPc12CC0NYEZepTbaRLph1m+XvMJ4xZA
BGdzOEZina59Tj9tcSP56VWH/Uv2tg5pLgdn2mdQi8NiW1xakddmTXcF1Guj5F7MDE8rxpNdV82G
TxUDJ099TfCg0wqa+x3WbEM5dDejYric2XCQH1UywrwhJXw0K5l+iVHlclixNxNbTDyg5JKc/JPY
/UDFfnen8XZDGsHsTiGD/ls5Z0QplY8gz8Sx8ImYewMdFXhkZ8A+Lz4IuWFiGvSbL8sml8zKMvkt
kTrGRkQKyOKpBekMIwTZ4JeUrIn+saYtI127mQzFsf8OjEwDegxS9EjI1Z+ZMdu3rb6L4VV0sS87
f2rzK2kyhTV1ah3rrOlO93X5UnkNgUM6eliuEB4geYlcSwxTO/i7+MbCU+imgLFwdKR/OV2N1WFO
P6x3iZ2OLMvjAb+NY1eJWGxVid3qCZYuu7zlvvhvDPNZG2OnpqSYcCth8mH73cSXs3opPDX7Xxfj
ks5DVEea7oQxsbrgFIwO+TUmTGfbOu9QlU7naEYom3kP+2P4PiUmiU1/bIivcuvFoUue9r0qmH6G
VmbkzKezglG+8iNarOGVakWkGf3e9xszsbgF/Sa66ceZKa9837EWd+XrUTrM1G6VQpCu89NIQ5Me
kU5zCGK1zLgplpUcud1yioUrZmY0cFfRWdgqUfEa/aT8fD+WjX9cRwMGiT/r9o0G2UdluUbS7y8p
xj4sWg5hHKvom9tWets+Z1Nf3L1kGRL/hbTfVGQ5WCgLSdL9avJjm00DlkuriiqNUA5XDvMeb961
YBRbkiv78Vv2kE3HNPl4g6Te5Arq0FiKST9h/rAFst0k6CZvRhNjULvkuIqVD6AC2wU3KcYEFW14
0lZ0RxHqdiojyzBikRCoMb36KLUxGYSpwUZue53K8dIRCN5fJxXjq7oiXoDhqZQ7ckTzaMnO6cTq
7RAu26c89nQcHVNoWvZU/IzKOCAJEyiQnLEBHWn5bHElJNHB4SgyewtqNiv6FIR9EIt2k++6NTjA
O0lzPnjVZfexASM1W2YAkNDXpLrqv985kMr7I79S/QJqnMjFr2lYXnTAV4eo+d8zZzj780UkoHrh
puVz4tkv8VDLqVW2vYrruLItkBPZ9OUTq1HMjELwc1K6FHbnlJKUg0swpu8+4icUqcygeijZMfQJ
JWQSrdYaVW3py/eiGTcxAkV46vM74V8uqoAVneth3jmiQN75aGFN5hlFDLfBXC3PNW52l3TvKbzf
GnRv7Mx2yWT0OGanY5GL9cCwbZTJ89mOWm97Wl7w93jfsIF65s4f+96Hv1CD72MC8yi7T7roCYYx
VdytaqU3H/LAsBLcYVlYzFEYS37G1glI8at6UMOJJ8H1b5bON4QAomWbD2o2QbOFlFaV7Jtw8FuQ
RCbJW0+XcZ0KaRieawI1fPGQ4XPxNahZ1Y8gP+NH6omSu+FGEGceUrfD6lXc/+AxhbvIqQ2zDQOh
xb9qIep9Bc7R4zaCHqcgTHVfdl9jXZgra91CXv7eIPlAJBuGBfdOSF7qbPJQJMZvgW6YdklqegZi
lL/+OXyZoZZ2h0ACAKRk0V/1aswgyD2bO39LzFGsiAR/ddo+LYqI3sEaqLoosvleRxzslN7etn+g
aacunElL3w2ruzvnsiQo/iuK7OWJqdSBgWYu+jdxtRO9N/nN6/Io4OXoJhcP7yKeBu9xXy4dhxxR
R+w7+BjtY8VM2uoR8PU8QYxImhg1NCqV+ylh5T/CR+5BP+KvfJQfLVh/6nx82lj0Sv0sDM6TYl/O
9Lf1RGe1KGSc1xetzvzJ0T7TJXzL01n6TxMiDxAMEUSw3LobBIcPC9XzpL+3M/eEGgI6EFgwilMg
fqPBJW0gFsegChk43ihK5Ltbuvvd8LpW+1VqNs3On8a3apAm9cczZiUxsDppD7iWpuw1L5BqoPLt
R0Jn0hib6Co9UILuivbjkghOZ9J3/mi5bZcNe8FOhL/Ux15Tzx88nSwWHIlFcR04n8NWp3bCe0pO
pmUHRVCyaOXcZFNW6hCsLRNkihFqyAZE4v9UP1nIYzGclqSC5SkVcmNGy20eqhUvmwg7x379tfCA
y2q+oV2W1MEPFtwhQ59kBrqNLxAKS9meA41Dhy+jM+FPJ2t7w0opbt45Gpo0wTFi1urAI6EuS/X0
oApmcmqb32LhAI1GLLzDGTH0MTmNZ8ArnZS8Lu+APa9bPxoUus6qjV/lTOZ4yXF9kZHtHx3Xc9en
5jmAcemfKof15Gln1MK8oxcZFf3MAF1L3CsU4iU+xdTm4azzpDjqqIMu3/Indb2a82Q1x/STIwwe
JPHbs8IGsA2/KPnEivfeQnFW0eG7JBN3+S6amowzn3dn36tjls6YCOiQwOXTZhhlKxdX8eM1ccq8
suwJ1hWQUstghIYseHlKVgixwfKvlCfqP8q53JC/DfKvRQsq8UDwa1pwqhFRbQNppSHuPrQl1j1r
npxsJ1kbLvRvKh4Tves4CCzfeBh+EvU+zz7/Qi4/nCK8NwrwwPOXRIYG+spheGxd8Vry8Dt2I1wM
4BF2jyAfbTPzW8vGzg3NK1A4pHwuW/wNJghRwPF+IsGr58ms7E/9cikvHFhRA/0+ZeIpQZ3BlFeh
7+wT4nb5+9nNWj1+ebon2X3xG/NqNCyCLNzaUtEP1LPA1Kol7k26Nod/GHfU9G9BkDshnft0cL7Z
3isxjViQ+IHnZRcYQ4CTpzpNpyYjgLqccXhu7JGPCNHqdch0xhHkStZQETK7s/pe6LDgDAk4/wDw
eVxaQLAIEhjrOxiB/r2oEAK7zG8agroSXn0C5RMIOCCVlhz8Iqsz4Ci2O69VH80TZzfDzNA8P14i
mHyHWEta5ecJ5MxvZ+aGdOmOYkOIuiQDLzDVTq5DlQZGezDSAd9HfmxMsoKALZFXIhiSK95J9FIr
h5MRD3M1z0Qxm1wZqR5I6IFNaqM29euFKidkE5Abm14uDMtQuvfCd20oI81PpGfXgZurvywZOGK9
RwKD0U6fUKsNz0FdLSqRoz9bSiUkN+M4vJtCchhW3bPVhbUQYc0espzDlVanmHrlHFhKgdLgtKai
TQ3MooviaG3jM+s3ommEkYoWknEitmySnlZCUQZ4//eIEhk1fY3ZHVfruhdOYNSUeNUkV1FwfpJ9
7Ghs+yfgEeO9zibcy2pQCdAbNbMYsLpyNPaB95Dsh6eWu4/d5mjC7lo23+OE1bVbE2O5yuOOzqCe
RzVXmSBgXcqYM2xlNK1bw5GUGvqjqbrfvA0J/svClCm3VZmWD5ZmvHtxJWc3cHNbHFgCzmvHeQYN
aur5yl7SpCW0kPQnq+dZmCCeA0MM6T+X7yFSKW1noyZ72wXF9ufsJniM2nTtRn6ujEBemG6uUESc
yYLzV2NM7JFCWsT2X/QO/5Y0IOmJ1k8TQelkS/hojx+DujXOV5cJQeKX+fan2UeSYlP2tvNZRg4h
gObQ7ewmUyvFVAHMGih1IVBQbzm/rVAAMglqyUR5NYgqTYiJv5slVLvP6sh+wO3RSATj3xlUl3uY
+RaxEAdQ1O4kuW31bJW70aOpuv91NmLqHG6AzkLTxdE8c182etzF7hud3zPkTa1Uygr/TndMLZ+Z
zVo9Vb1QNDippByKs+F07bBj9KKy7IjDhLhqpsVorMX/1jf3yqKRH12VqtVbbPqkxXzzRSbfaQ+W
R8k6H0bW7cl/Eo7Huxt1uLpbglZfUQE2PjiaQZhGrQ6lBTcSJoFhcAQ/funTPnaOB8LI3+d2GB1B
P/MaYM0Hd0CV/kLWO1gXMB7yI6xUM4Mtn4bEhX4nbKKAfcA8w8eu3V2G9dNtBsp73teiIqGTRO8v
sq6Q3YCO+l1MbjRiycvZMmlaUhHon4PfErv8OGKb/M3qrhUnqSnLsUAndG2iZfv/MLDwjmCGJQyq
SqSlWA9xAiZHzAnPTM28R/wQ/onxzlpLCbC9/BT6c/Se0JnFci5ksIxSwcG/3rUYsksRHwkT3cXL
M+ph1zbOs5pzD/ynKQryyP8cKqcp9L+YuMrcHfO2GeCWu6lQUsiIy8TEczlzZfMLlJdY2AjRjSKW
dXCYAsBGXupXfvrDgV1ZisZbYf+f60y0wpv+rUgK3rWO95vf29VNDe+K1v6CabQpPw885KDYaFB0
xzAL2hyv54hlzHJ7pQgmNpiCX7dW4tJT3+7c20xcWVVT8tqpQ9u7VcnKB/+NFiidesGT3oLpAgwX
vfXNQL6J+F6gGXx/rq48ffqRSQ3huwb2ySC5ASQ8JQHlTVPg1ECXbDFqJL9UHpBCT2eEpNr759gU
Cr2+st226MKbfmBnwEy2AWhoaf7CL/kUKSb5I0qujH95qjDqjzebIVQ7aslPzFTjXqXnSyGwAbO4
tkFZp+BV5REf1IJ/qpnGaNyk/5sH3x14dozfvj2xmt0epCiDpTVaNpAAP9/koTa2j/OKVc/6Tfhz
FICctuTP8JF05TkxqeF3DmM+6mo7k6spr+B4MFxmpHfi4ljlpuP1bnaYbb+hi4eWvF5zncnZxeKP
Za3FWMcoe0RvACZPJNvFhYdBBRw+H5KQ+54qJLrm8j99kN1boN8fqb/1cJTU0MIfubqzk+mGUAb3
XQ3eDDjTP1dtKbjmVgbxfKn1Gj6+Z0aVewwulQ5ArdVO5oVW+5d2WObV5ItsABX7JFCHmfexYgAS
erepLRMfIOtWvKPSh/4SfJicnnFGBN7ThkhAQNnePyJGUSGk9T80GePpM1Wyf7QNAfFNltMRbR07
tQwaDbhkHjgsvLLF9N/cA6jxN5f3+UIgHjlTSIqgEFVWqQXzDiiub++jpF5tHgpCqBLuwUwuxJTD
hzdYFZo5czASO5027BTsHLbtYNRak/3YpRJKugr2orKbaKKXlkkmAHdU1k7TkFatVt8dGfDZHgug
4lt1JVaopQNiZEYkAxA8d4DmDekgYMuzKR/9y9rztlCJ3sEpqXecD0ExcvLYxDgfPVe3N3zMQu9X
slwvUI42anXfU7VmvvUEGvMEUIC7CuSMwgPtKUihD9+3PCCjWmr8GRr+rkUHuKt/TPJBFe8qhaNJ
bDZ4LiSzqk5UR3LCM/1u29pxft+UH+Tw9rq6LtgJLE/4t1YCUSeSw4M+3XnTYwqWyCwHdYNvN4sc
A0wmgzHH/6Vd3whWZ6lRJYNO9H1RVWQVG9Qqic1k/6I0R+0GBVcVS6Co0VGe8PzGFKLIUaoBpUZr
k0bcg8nlcBLJzTOxhEwkB44h24EocWM0H2YmghjxN1GhI8p0nasEsKWiaHcPhjnoVnlLvVahWWcP
ap3mOGJqJAwU2aXP8pYy5O4dDZ6uhyJpLJHCKO65bICAmyZkaOjXfjbfvOedCyBho3FTL5HYt07L
8Krd0aEdNlpyUVxrR4mH+G5AOsJ0+8vacYOvS5Q2Y8uI/QjUjbOx47H2TpzupZgRMXRhTfwAQYmQ
oeyQnXIkdkE72z615sE2ACH3UgbnYMMEBCmWZ9b6FRM5pTW4EIsMb1TdkZJRMz7nKydBigjIklPY
lXgMAPXQwqqDBAHUv1ansGuB23WbdxkPVuI3/iOr1tqYW5g0hWbMK8Bh0JFg0eCOd+8TyemKJZwY
e78Ue5UPbURgYNlpUmv+uCn+i1OUoEL/7XD8BFNd5jf7kXNfzfG+fQqMKjXRcj8T4NQ8GDtdPxmn
xrOHYzy77rfYSbklt4G3N52PxS9ZdcWu+jo/TcyaeO14GS6hhMuQPHhj25cpz6cHTvOwFAvzQIfY
OBHNm8fjz+1+t+08VB9dqvtsOJPfFJuYBjAWNCDPtBraD/MAiwdIPTP9z0YGbfxSeRMgHilShsvH
q7w5uQucF9eFGcTIssqsyF3qYWGpaTRL0TKVU+HclvJywhxVSdSYh7RTKF/A3STG2MnXRH6KCDiE
/mYflMxhM73cUGDvhPYBRGJk4513M5ZrMEQ5ymASjNnbq3PBNG+XF1+7J0szoJfa7UfWaIaVi8ky
WZnuNu3x9e1QCFfOMjpe4dPGN4+4vIjOMT4A53ADgt5tJycitdKgJgPIRkRv5ijE3cJFIrDoYsbA
or2c/4jkxSkEfOsYv1gD7ypGm5TvghK7N+kn50lmHuQIQ8r2oxbeXAv+P5g0RndAFGi+k1XImvIc
quGSs08rFPeFTmaDF9Ue7K/YPH0xYY01DfxeaqAjkHg5wAEATNgJecrPYUBPqnOipwsBxUaleFSe
ojkEWPGa2Rtt+NGN4qf4tfE6msNYm/86YWDpoj7NqKrwTbeVOB2BjdHtr++KwnnE2+TW3h+kGpjU
A0OiWQCbKAMAPxE61dX728xRWRYYYFu5yZO6xJoRrXQvaW/Xs5UzxFt4ZGib8a/wtzTb8jru1oKf
DocgLH2CJLwXfWPw8/GVc6u4VvotxwRkGM115TYpGHJd521HKXj227hey7hjRgQrnOBf452MUkq/
OtF6PKA7T48NEJbX5pyebnjcZvNRBi0TPzy3Dxx+oxvsH6rSWEZIjoa+1W3wpYfZnD8s7ns3i8mL
XTGu2YX7AaDsXnGd10Jw29JgrP65Q1ksJfWKS9JI8bokltTWvAxBVwh7FIrFdHLYIoqyJU877wS9
s4ibn3FnBHSirRHjxDa+GVaDPNBztufa3YfFe8ahDZbqUV0cmlRODx3eZZmT8iTiOlBGqFiI20Ii
JqptpG0OLs/i2qwU1XalkveetsbZGS73upRwJTH4pOSTnS9o2uzz+cFSWSFBDRh46gg7ZZNaByo7
uDuXSZYSIQRgZlhS3pbcl0Jscpg16iqI6ldLvVfeLQkXP4x5wtHjFDfC7liSKp+1WB/9Z/WkIxbL
CIFN7CmI6m0eNRBUjgJs1CMOBfelMdfmReOcWrN/Y79p1AuehA7lPWl+0bY+0rTAz/ctuGuNY5H7
6V+b1yF7smW+gqGoYjBafwMF/pnXy6uNRo8h4FMcIoluLYs068j8gqK7rOMJSJ9zCNuIDq2S1/Op
8tNg/jG2ieM9RZJKrY3znmCY3PB3IUilakv/XZmAby2QjcSg1d0rPH55UUycRKOUcE+8tuijmoyC
WuNP4aZu2AP9EaQgjuXNA+/LGW/rmfqJy0L18hquppv4TeFjLtlniqdcaZahW4a8VoRskYfqd2/b
9OoYvJYbH8Dgrppo/p/vOwlgidZMD6YDHnKTs+J3pkLQRhkQPdHto7pdMY1r+Ks5AXwQ6N5UoAAf
60EO2ZrlBFWmJTpzV2QkG9oaCMVAkVgPZWkO8cJq5J31D8Dqpzj4RZeJ3fWDyJUbL3/o2n/nhWne
rtqr9o+nj3IAG02dcCkQbNwizpBISVIGqwFqhf8chGUA0b5Tzl0pm/hFjMrFSulFLxuoT+xL3HIK
sDxOii03JmFnCH2C48s6fAJ6ZUQuIKWHpWBbYBRxixyeJt7ed6/BukTYicoNIAhYyuKqBCBCGJtn
HbwI+qEhVYCS7KJYO9vxQ/7KkDVvfqkWE1xMm7zNdgmpPiiv9AKiyvPlbETCvz2pz9KyyfK5gy92
v9CiwXXk3UDhGdA7WB+NTp7oagn8ZzkTb9+Q13ZniCIMhtsoFoSHgFvyrpddX3cv5cUGtzShYMfd
HqPTe4on3gVIR50jq06HWtNYFhZXGpTP1j/LRAUlpgap3cncBNhKaNxz+bZnvdzvSOQGfxcsoKpY
fJBnQQY3/O5cYjlmdKcu4cfAdKLLnEWJEFBPNBByw9f7uEKacnh7B9+GgdmHpDnvoCo2XBaRTkpq
aoiagn7PA6097B4+IwY97I8vCH0BPHFUh5fOXesDd9S7ZbDPrn9lmXUWFzGSG+evPbfa0oJgm6qd
NLsZy/rcUv0VAgkiQaRsj0pjTpWWTbHA/AhTEfVJby8JHCvYm/puapVPzpUgkHAyIbKWLn+LRFT5
VeU3uG7ar9AhAygi6lAt8l634unIhJmhaR/kItClEQ95r/iyCCEpYqRDrOkxDQidCBEybhx+mXUF
tarMy2ZgXxXPhx/lAjDiMdF82qLTlcKka1Xc26YhGh62iz65dw9qR0XXFcgXYfXqhoUy7t0bKs//
hfYGzZmzsIdhHSn0nvVLhjzoK4AKK/20xREgHX6WTS1uDbLCSSf2gFtHiW0Y9vs2uXUnlYOkTpVX
8f0502WfVTl95s94JjRK7+FOL49oGpXdO8oUZClJlAUDEh8zYw28VPBI6aICSQ/lD3ywWwpEC54X
jc5jQcBrwb7PbcwgXp10Q+um/CAyh9Kl4hBImPs8UbQO82c17bjJqAL4khfS5+BpxI6ss0trJW+l
QVIpa658VuGsuU8G6I0Sh/lTu+2rSRHJXc6txne6MdH8ZvkCSt3x1TceYfHva9Pmmah9M5QhBHKd
EndjOo7HYpJ+qD6TGjOrIAcNfPONxR0mLY96If7lD7NRoqa5ppCsUBcTEIACqfPhavy2bovnzCkn
P2moPTE527nGxck7LrmHxA4e+nltJR/yAzqFeGfflOkHxwzJ1J7HN8H/Mx09Y22JazpIaP2qFR2J
Nfe9pk2wwUMnbQTqwEvdoQLzCyo3FQStFmGp0PykUmNbu3P/xt35fp7LEBZrDstDzm75QCyIi4bH
it0D4GgOp6lIUAiYtKkFyVv9zVgQRohIrDdLJ3WZ0qBllfi7jTjsbTgLcUdtxhtGM2wF+IY15HWI
VhSPqg0mTb99h7fI/adFA1aWIaTqGsa2EmKL7g84Ul8xwYPMbBL+Pk+83hrKhWghxO37PN0B+c2p
uCGLC3nr7ACo/0qJdtSm/XyZVaAhDbQl/gAcSnCGRyiANFgWJIsqb5lcQBELAm/n+3yPY7QZELxm
L8wPaMQ+pcE5GXD1RWuqNFQm2ZVKoee5xZzr5qlmlwocQAHLEvmBp8P042MUUoR5OqpPdjuI4HAb
vd14wrA5hO4iOKvYgKdFbsG1ofzr3jPKuCiRwNzh71FUQPEKK26q8cwQ3N+Iy86WLzQ6U6OK/fd3
sWDzKQ4mB22AeVe1+16J8sqMN3XeiJ45uv2L8sT3QpKMLlW+pdPrElOzniPP7SceX6pYM2xfYemd
kwsAUX3iZBIJbrHi7kef+eFgglve6knuwUpCBB+8lSrkIWOp00oaqJLlZBI0OsT5t3SlVA7E6dn+
7Vg+iLDeoSZoqgb6APq+7c+NV8QN2TPcjsmmosYk2RZU3p6tMfBfBGhxr/D3wdLRFV42mSw1U8Uo
QQ6D67ylhp+AbGOn8hTHqn5x13tbeqNJsoxk9h/JZE6yvpvqavnzpw14zSVL7BW+8vZobpLQdxNw
Z7vuYOuEILPX/NEUoZPirvnNHuTxYYx7Aw6O3+02+k42n5CXTKOjVbQ2JF2s/2GGDtkJRUELACiW
U0+pz3sxZZnjiNTb3wqAAQ9X+IgQs/xwIRynw0Bci+nS8O4zRodn/u5HdqZw7MLubesCpgzL7UtR
Ic5P6KDsBifxWY2UGnI/QgNTn8bYEA/zUxykrKVdfE5S/QiWa+rdHzBDEv8CTPSsFuANhPpW3Ywo
DogiXtd1EJ/D/UsWB0ESvXfCs83q2vSGD7w0GITDwNWIoAXLYAODg4CrgzcZrm4MZlzUKRRAtTOq
9qJfYPsZnouJTaqeOzhyySiVPoxZkuho2W/4sAtFvhLJ4OnxjuXyoNoan3vnT5KYESQCO1Gnhtac
mS937wAW5+6IdPnEgnq4Daoq79JiRiGoGrl6GL/eEoeTQarbWuLXwnWnoQApmS9RQ8FVc5v6ZtKJ
6wI0asszTRAEkIrzuuM4xQ4sy6Joo5pB0zAXJEGKQcWa9xImyq3oPUq9W/DwH+SWaZwmidoByNu6
9Ey7dUwVcvV/ki4oEKWF7fuBVYSS3FFMjveCYdlanE16QGeptRhET0cFvkIqR/wWoNAsuklPHYsX
WKkfXZiNyvt/xfszEPu1qMldosiw60DWpoMwI0vCr2CEmJUq0PRCDirbdVDu994pQT3ScNd7WZoq
m1tRRaxER4Kpz04weXhGe2unI5DIg4tKsO8uHWhIwhyRfDOZ9kat5mpA8/HiFnZ+gfHzfaqbdX/B
VxWVFmvNAGCr5RyDqIKQmkwtTYMV+ZmcrXx8++Frq7ou0NkAtmNnNEbFMd3r7x6dYmKpfW2/68oR
fOkWsKShfexn8hiXCZH3Y3cGu30nrj1Tr7hRyoi7K273icY6aXOk9BEcOtg+jHXmIRf+OS5QfzaV
EPPJeitUWHLUSjA/fOwnCiT3mGJSHRmp5YRPijfft0h3RF8bXN4jLaEqY3hlR5ekQzw8a4DUvXGn
15cRBKIPw3O4DBJM2+NAuBibSbh3NHGWWK3UZr6b2XVxb2rswlf/kKeE9AWyNnukuwRaDLmlCQ+J
R6wk6C5JkV1IDIM0RJUGPJHGK3EJog71k+e8jLs8nCLocqnh8V8Z5H7idGVlKG5OgtTKYtlcQvZC
AuWY/TxKRONDLhkCa1r3pbmLJG80pIubDjUYw76FtKM52bkpSIVljbF5QpWH+wnuu+4DQANfsXtf
Aq3CEYesHsePjQU30qH4YnPsNEEhqOXv2YMoAf5QZuBrLIfzCkfp9DzXDLVyIMZnIiVLd7w2n16w
E/mMG3QWygC96VXiQaYBuChvSowXx9pkkzUt/UBNgKLTrGT7ZEHBw/f9JgijEqd2EeYwewGX/Q0p
BWU+QQ4Z0rxRejXxwwcOWE1QLZ+uZWIDjQKD6mtAZ77yDiq9aBYdd983yI+o7V4VtyBGnHZBu5QS
euDeShNJkB1dp2QibkR3NGq+WeV8AGxfj8J2y0c5IwwB9r/uJiMaN6sqNLbHNxn+N79Y5Bqw5yhK
3QJKsW7cr6bUwF9dibL9pX95Xqs5PlwDBMhKJ/fmQ2viIMDazRXDi+fwqi/yIm2QMaD+GAkK0fsq
CTqEV6z10Sx+ddP5jR4oc1xUP15c1sUZRpGXQfHbA36HyCpRjHt0xC3bW3kmHVvssIWEglfPl9q/
05/uK07NTiQsTjFvtyIcQsOBQme1Czd147AD7m42Kf1wUwcS9PwOkVJX+Tz+kJh1wDqOsBAZP/cA
DnicZtva8TpOjKkb6BYSnhQ1n1Na3WJJnouV4/KzDZ/7Z6lKfiet5e6db3Pq/zogi/3p+4RwPKUV
ues6urj8jPXeuPVfy5JVinAlgsmZHhG+Py9eWmjF/eKS0eLhImvDNQZ37BL301vyuAV01YlboC7o
B3Bc3KxxbynB58Rynu4n3IYKjN+sYgX9FyAIJ1/iGr2lKGn/duXUfSz6rFjsI6T+DmA1C8gGjkIi
DlNAVQbLE4Bge1rWTv5/VVEBIUwZywQ1m8UFCymw/ThmR4wqyU+k5HT8+C+1EaUQKhru0G1DpwzX
DoclPYFVQ8hgnBbDkDEkXOlWEi5RKCrHEJ9HZliaM69P2ix1HaJ208+KaxYFmMvNsxYIc0uvuFE2
jI0PjCukZ+VnRsbRBQN6QWhyAomJ8bkWLhRr/8BUUiwlmPwG/ScDoiCesBe1JIBzOnHq8wh0VkwA
CN47tYMZqRH/evTrFDtgMfBXtOi0IHwcLsOAo55U9mXial3S2pKs9pNIFMzH3dK8o2b0oGr4pE12
6vH5vJ6Cdn9xXwVDNzXe/77MeS56a0GmywdiqRqaDQYOLST2zHFEyVbfFZe/iQXyxTUBHtuG1VWO
JFm4F5LO3bn5Mv2LdJpMSw2xj5CwbXpDt7y50qxB+Pu7ePgy5WNsqURyGYHjtFcCVwPSlYPvW9F/
nT7ZHi4jpTjSnaWwZmxCAh6bMnIrshq9uzUn38adkPmyQs0Y2gA1vCCW6bBYZyHKhobzdrfrrJKr
udcHjvWOq8EGt9HhZi+ANnr5ORs7tyWEcqbRIRhdsA/kBVUC1OtvjzCv8nGW+9aHnLbE7rkCLD9t
d27b8fsruXW8nM2u+TixrLBeR1+R0zEMcX1GzTJHJXm7+XTNWDDH3n9d5bMRpALk9SGdiZ1/F2rn
jTnC3cBvphyJklIzeaJ1o/LMVRda5q8IwxJRS/zW0RRKl+H+IJkH6YHPKUaCbX357o1z6dVisRyO
n01vrU4plGimmt0lmBqixOzZnS7t6Bdh0+29R4XiY21ltQdYccM2qRUcanuLparTYVc4iWMqy0Bg
0umYbvisKtYtRpfiyy4xSN7c/LiEjMkh2rYCjmT6eS1a+0Eh96KgydL/DtpaDyKEybks97VH7dKt
wD+WT5BHaAL8/MP/0u2NkomuANHWTu9BuSDV7ZkbC99WlJ9Euyv53MW4GSQmmg0necCWxOYOfnvc
YWdcYAaaVQUr/6EXfSgDccGJHIQFOyGD4baA6q50mME//0ghjTDIKHYHSDE4RWCZ7taUqN8qv7ME
90Qok9j1s1LhbLCfHKTx4HamOGq6Re3mb8PBfzIBPGOUeXC9Vo+rfitBKnwhlOszfV5ox5+Y6Lys
RoZtE2Xy7Ug65nitICWmqvAzLLdGEwlMipAEDWAm1qDDWKsr+uUSmTwW2JQ4M0VZkLukELcreAK6
r8H1lxjwczu5RHbX6Bg7wyNgRpqkiCWWD/nBJx0nzBl+2EdMNBpoFnb8es6Suwcp5uNtOxCPRxGA
+zRapbiTXbcs1Yc5UqIGS2S22odzI0xx6JcGay50yjx/WKJrYgyoyo2J1u1l92ZfjHNMLeCBrMjM
o+Yt+Wh6P4wWsHpuC1wgcCBIzJN3Z5zhR4jVaBDuPRA/mJ8LzRmsvVnc4EoEoTPCDH9fm3FnoMYt
s2oVnvbuzNjXOdo4AnOikbNLT7wNJHR1o4RtFziV0LI0h+MxcFUun1O7iCyFc64hKHq4YG4lNF4x
miBfZ/wTPtTlWgzT6orJa6+kK8FTttu7OoqO0wmJgaopLMo1W5PSDpJWbbJpSLb8YdY4QAm5EDiN
svpxqSWzA9caG/sDBMACbxjWzLGI53tc4dymozmio9gJl8Y2qsc4RMNbJpK8vyfmL/CZiTA4bfuG
GScwCqQO6O+by2Etd1JMf3hIOhiu0D4TclnSXj5sYO9QGBEAxeJEhq/2woFJJRlsfZsdwb1HYhdy
E31QD/Xxh8+Rufa5JLbLUVj1QVlsQkdgjJXPepm3y/ytZ6LEeTThUucD5ITDTelEjZZ6kWpSg8VZ
NtbyGKRl3abnFM5EUFxn48+G7hZwpETyKT5Ma2DwnDS09jtAi5qOL0nxkl+NJozY/pFWtpTepbK/
QvW05ddf1oSNudG29rpYd67DLN0WWQdVv2LaVcRtgzZANQ7Idak5/afMVPf6xaVK5F8jkMTfgj/x
IOZDGiwcAer5feqNL2FiGEx1l2UhUlNiqEjMSXiq8xj8mxcGO+RNosTmxFhffrjVPm9AC6g2eZDY
hcyuHH8i1z1/6kDRsN+1kpQSVdu18CryJPlFm1Vq/VZY6Dl8gsRhXlSttvsKcR57P/n9WZxJOdh7
4NHxRSTrNOXgtntho7gVRUOlKrUfNBkh1WJMxiQQxHBATusUwRexxwh0HoP3Rempzysvgd67GzrU
fROeY8ve0hjB2YuHfxTWNuPWuMlGmyXgptT/FBmknOQfX9GFKdbdcZpU6xRFYrk2KEm1P0qcfFdj
B5MVva7q5XWNyFf9t43xNh6QiXsXrocjx40icIDdFT5E0jxAmCejXQgHD6DE+eBc3iFrJvssdwGn
t/7kUFIuGr3ZRQZeu0EJpJAf+tXFlZQtbtKjmfwX1HRgrcnRoIBzP8wN7ANnVzixCPF8t8xCRfND
/6w/NDJtm4u2W3OsbhtAjARYr7epkrNTxYuCrJMAm8CMY5wJOgAVxHWw8mm5JjYnF0m3yJOY6GdW
mEmxHu26PixmTURrZfkkju5Hrj8jxAy/K/q4UribIqBr40Qs8RHdstviADohdU1LxZ7pWZGoSu/n
nkcJbAPPVeONj9mc7+pU8VdKr494BeKZYJu2s+YaHRN4cCxGZ0NC/V2jnrtkoKB8BlQw0G08Jm1T
dD2yRVmcN7Yoxpuku9faeZy7NQpQ3nbPai+DMDxiEp6/YIoIr9uGQyZOpH2OS44Dfljat7Q3V17j
peRf50Jgm//mEBYdNaMhj3j/ictuQ04E3QqBaCmKovzYZzQd3SujZFIF2nCauRknoEOjLND8cbmJ
v+VLdZAkxs/5/JcXk2blOPghf9MG39RUjfpzaWdtTZ2VeYSr/5wBNpEz7DO4x4WhYU5+oLbky7b3
zJ3du/mlu0L2QQtU/0UfPFa5/PyxGuw2rFSQddV8uGG05cOuvve8+cbofy4fY8lRuxKTfEMmtsDm
EtQBZs/FvPj/E7TPRqUORA5OUigebRGdW4g3P7p56qLTgQMjexc3A0Y7GgZnWYPxi/I1Rrfa1i8w
pYou1jGug55QTOMX7ejITAFXM4UXpQPrIUSwdZraVoNQEJ7l/IJb4ZLz79lNhk/TNR0Y9faa2ZuQ
rTvmJl7/UdRSmUwbceIqstXRqGscauQ3YmhfilJcY5oylnNAymVPbLUsxsHTOUv8nd8/eiVbAvqS
Mk9loD4F0LA459p9JpcxyE9WW+56He72QsoYWnE5zceR4LKzai3jvJ5XKLIL8yigkPi0EMkWwq2D
8hnALDJXjRHLUvGBUv5CL3nq0qwxOBm0cUVHsYDglErwGJhmdxgbKZvTe2aRdqQa6n3i4pkCwS+q
72SuoVJahsMF/0XOSlFTE+6q9SCRxgogCgAazq2ROO3f5W4y0SgwTELnONs+JEL5hBf5asZYx8QX
oIQyVg3yDvV0MEVUCD5a5c+37Wjrtlrr9eawsYzf/mn11AzzZr2XNln7JUlb8kDZrBp664I+n+AH
jNvTNNPK6FjMwqfVCs0Sp/epoiDYZq4TPpKJ7qP9w1X8T6vMtIH5jXhWx7wzfzzA8FbkL0ZtqXrT
+zwDoajCF9oKneZl0i8mWreT4DuzPYUmz9NWoJgcftuXjidR/p2/EZrvVqOk4zaW0XB/AjPpsaYL
MWenT5+FOvHyBsoQgJoQQwUzJ4uTy3ZAS0XsFXUJZKrVd5zzkR0eQzb1W8VkO/DOL+FVvpvRlWNX
U1ZHhPBIf9AGan+etS7icg4XGceFDUv3oSm5m10XCk5+Z910SnUJvCDaHrpVBrglyqtnE421iqEv
yLInBrHhnL8S33ki03XdPQ4UC9Fo5Uz3WOOBDUal+oTXCKLS84L6TwoB7mtkBNschZV8ZnKeYR6Z
O1S0cmJao/4EWxDhy3QqsWTm3n9Syehk6WOsU6SUxBOoTNhfeQFOViUzO2vIGYpNi8jhRtGZJ6uc
CBBdswU43yDammFLRpWn50UVRgF0aEjR7LNhisIg/hCtTIkuVX/pI+kyUmAKYBE12RhgL3pTtWw8
qdZUN74/MjyD8aUIhvbIalZGbawU83Bl9TEtUXm3jtiR8SvQ3QFX6xUUa17jTgoc70TO8q6nYT1+
nunhK4QFvIfGwQZTFXe/iybr/DEi0v+DyrB1V1ytVYnzlRxUJb0sSIZd4qjK0X5TEDp1Q9KwhWjg
DIOnJsZYZBtNsWAg9RESrW0PyoyPboJMMDbG5hyNGCDfwm0dC6OE1WnALGk90gPOcr/j+tR1zAmR
MFDxAxAVI5vw7qGCinMA9MJ62vBMw8ucV+TQgSNlutKdsO8OANrDHhz40EIAbZhf8vTek8YOujfV
oFe4C9tMYLRK0+3mugfUTWsLS9coR7YpzyTbptJjJRELUrCRi6JPW0mT0P6P/yDuMcgZ+uvkAyXK
EUfAds8KfvrIg/L1oY9vOEd+RPbVLBkfKliPIqDig4EciC9l+NxuZY1eOQwqMJb1NkgacJPGBaBI
hDxxF1jnb5PGQ1rgHGrC52gd2dgxf0FJISm4gV9HAMR5dc/7z0qGLj7ta68oM1ssTSxu7YwEmtnR
ldAWk8EVTw3jZt+SFc0P3E+6UhR2C8vFmlqIeMLnXeoJ1cVOWXBwLPOvOm7ojd/4t8O0zIROyHOi
pON2NFIE5skqwGWLdNKZHQcGyGbeiLXwOTV4q7oCAiENT0aaR9UYmVnLMm+AwOYSeHFaN3y4G5Qk
AJ/EpHPnZCOTtZ+kCdBdU2cH2NM/VdZN3/ymhzHMpin2PnmjH0wdvwR9MG45oMSzoPGeyyxtSt4+
d+wjstgDg/raYBbEPPwPypPRQ4w/OoHELVdbnOvHGJ/fOti1eD/lXlRWtbsvP7R8jkZbm2cHnlEz
ayQT0TwZd3BBoC4N2k/Kz2b1Y8YCEgxGIX1su7G/oYjuzkV1DL4aitibds6s+34saTxaIyJ9zLYt
rMCOoPoFd30Z9LtkbjxDgHYc3Kt8aWG5TdO7J11ctJg7DmO7mdIUBlADd3bRi6pqIuVpLrldSt9E
8QuuBuHLFZ7VxA3EJmNCXU0RpfdFAzDod8ICl23QalJns8lwCKHkGysMhGKkLfFWQSQEd0aB5NZ5
DMBUPOXZIoq9NtrJ0AJ+jtCp5Nb1oWPZHNJRCCrpKfTUJzXMnt13mXmZhp5XwP7614c7QeiYTnQW
vhnFLYceumSk7uFWltF9KbvcDaT3HQS4xVnOglRkui368X4puY6rAAeWCjn5mNmjUZKVAX9itBaP
vpvmUmBZmxfG5xT5TmVDGfAGa0cA6zXKZU3bRSmNDRtvWCuCsu5wTXrbR3Hqm2y8DpxXnVknsG3B
dlM85SMs4NXVI0z9VRKjwM9LtBBwtp8BdZ27Lg7eveBsDXB5LSvolYaDtP/CuPwakJ4GNQWiiSIQ
eBALkC9SXFc9L55K/vUPYIKS4Mx8aa+/A9xUxzVpYzwIO+9oBQhg6pSM0y3KiaDUcsoYd3gKsJV8
YaJOTVtzhmn3YRbH79lcMKrZOoepVuNJLNnkRaN9CWva5nTPidd7aIfOK9Tjvm5ByFirjxTeNPzD
vTR9CVUsygYyM/8MAcERC6B5WhQPzHzZG7Zn59eyIL2JVdsEWsLFsapsJaxcrKd6VmMFT3M1zZRr
/lzmm+n5aYS/MLL204ngnKbL2pvi/+VYdFLKYhbB9L1Y8U839ir2FBz1gNYzT0bos61rDOTIo7pR
uUiI7/v3hugClNTseHiYn1cJGJbjK0ey3iZuRzMjXVpRplVhJgxu5xDX8q2Gl1GNfzkVSrTqVUax
+PSPPuyUagnqq3M4Q60rLu1m0Nmk08sx4JHwekqytfVnMQN2cQ1shZ6PtFM9/dKUtGLB4MFXVCv+
97cS5jYuyKzqZMHm4aQBDjDZLl925NngG/egY75H8g5XKAWHywipRPr5IE1f3tCpvf/pnUyFoT6H
Gii/mIkrOMBFjFRzqroJjtlj46yAIISSi1yotcyZ9rfvOUgQEYVdAAvZOD4nWrpMrcvlctfkd4Q+
rOQNjDLRG5UnfI5G8nZAUvfWfDL0Rn6WDjDGKtwVD8/PEppndPuHNQVygsSUZiwNeExF1m8qCUI3
Jq1pR2/JDGiSoM5xUcXZQxhX9MbwIHFXRaeYAoCBxvi43Xj+R9brNHFYyXd2f4iljAy/CjNBLrPh
uE4gRRypH8XB+ygBDN+ITycbZZ+sgEEIzJ0mgzDJTltcOS0DK6BtuOgq4h5nELXAANaI920fHnZW
QqNanJh1GA4SlFyPBg9ro2kgAJBo9kRkY0VHS7zlhwkR5FppQMrP8bMioMld3VAyZnM8MrD+CVNn
lCJAeEfs5MMSp9vutArhXqDO2QyoWHMVgJG28N1WRw9FbbFyz1gowkHYTI0B8oT2DMjEe6pP1Gye
xzEtHA8pxlmoXQMrq1zUNusxq6nMGSpsFDSmt/qs6RmsQsdgYpA6HjGX3pgwS/hT+PGFmh3ie7Sj
0YFKdkyGc0uSsafOPEcPUm4TTnY4Dmjo8+82YdWLsCrgJF6G48UQkuRQfQA++RfYPKyd5KzPQa0V
qbbzZgP4jW3dND71CHBXkr7Uq7rvpX0+f5Hc1wsRhAsx5aTXCMZ3v6iE9koguoNwhTsdQBPAptCX
Tqjc2CLWh4+2TcsNZ9S0F0+JPAHxEpButq9zGNy9KQpjYPMOIbcoJKrjmWWb749yU4PGOu2lDFqy
KgkogPz3h3irkrZvkTVTXIj3TBwzwiROG78aYZ1W1gdcfDgGzi5pqGVb+Of9Yed9BCmHzPK8g5qF
6EHd/zYuCS3SE0IcfHMVvmOpw1nrA9RpnuLac01BBq/n+11WdjTiXEzuVeVDrLWTyhoJMXUUwf93
Xm+DdetrJAYfdgbtn3sLsumkYb4/78B/jAJwzSTPSl+tCgRK1oO6A8zutf9oWtW6VtmSLwfyBiFH
SJAZbZce7QPUkdvSTo1EJUq2gJAE8CZkSmhA6FPoh7N/4u4DnyOPqL5FjtFzIj9p9iJKMQItACFG
atw5i1bF940vhO/xdhjaXzYNtD5OZGLxiwnyEm9/wpMr+li7Ry5SpEN8rIhsACFhFmhlGwyPSR1N
kJFBnseIHthVXS5qvb4moadZEOtN7CfOzpWQGTj/JAkMOft9gnqdAK1YcdjOgAvPy4YQl1kkpGhe
YnjpzRLkk5egVIydUf78ZFedWwZaKQ9hHO5z4Ixqzr5hmUnIBIgwjvFBpFo84iP4PQcaERzVqFq+
tz9qbGNqR96zKcpx306R7QFh+WfHftiOruHxJMk5SaBiW1iSOYB3A8/1L122A9DB+TSYX7GKEn5O
Xxrozzsk1o5BsY8wWNq/iP3ECcoHvDZABIDU5zsfP+d3SV8Su4D7jN4NzUVkOSF1qYwKrza793zY
YOlNnWrlInr28/gDeJ0W7UuaDw1ol3tg9Otg2Oq6VudqlYf9l+TqeXpjd9vh+KC4PNLygxrHVJ84
D2FrdE+kVWGTMNWm/u9wtjGv1Ckv5pFVPgrXfzKXxXEG5YsGb7Xgwjn84W/fHA8idWbk6yvVaZZP
/pIUsMmA0PguRpbbveRTBZ34GMae8u+R04w5288+Kj7MFYFRbYeI7Fyc5Q4rJjx/64InENMFlN0a
02JWI/Kd0g3T/YxCGQWqR0kGIxrjV4p8UDxDW0fBIpXQ4NWlQKMHbCumh3c9Npt2icA/1pWDZhVB
4T68xnHgCCGDLab+1MWtIhT8TO5yBnC2FYfT7uzXVDEMFKRsmiDFA6cBSgaiWRxgcRFHNe6k5hCq
XiPnnIdvFlnbc0JfF1xb6mwF23hV28ee5/L8qKZkmXGI0Zih5OqXt5QExqdj46KnXPqpmHFnCHY4
eIY3tbr8K9NEn/dIbKP2g5U4FOHXy7xLGwZzU3pifyannJToCNwbtazl+xQ3d3U1o9Gh3pIvzX3W
9ZMxWwFPeKn0ekOZzFPF+T40txj0c9t3+LpnH93CEdAjMoLwfPxkPrlZnjKA8fJSj7JcLMrfpi/q
aAIDVUkfvC681hlmifYZBqurWYxB763r7Qs7mN65L2gOL2vPirVt3bBZ9kFYLikDuYsRhsa2LU3s
/1CdBzkUHML+KFKK/5kJ8dO1n3av94sPRNZJcrc60NrhzKOaogOAjNh6fz+dgL10fRw2QGMdbRad
9HlXItfacAOpnmdO6tl+f/UmxdVyJBcKwnhkHOL3grILCkD8kgSXVNzflE9XPbhFxU+TdQcbrTxs
qnH7tHCVtYuUdTzb/S3R90pBa106itRNIdFMg8eXVGvuF6SUvQH4QfA0QLZT5/3Oy6X1DhUUX+GW
3yt3LGeUD08ErNKJyxgxv65B6VQE+gAEAzz8Mbog1OJHOdKMf3tqJ1WjbyH+bCwOKBeF8XpXjhbx
f3ZnmWsxmC54qUTZS8ASxzQQn/RRwulwFYyTaO2r2o+n4iUCAzvRVkqE2o8SnvG304dIgYX04E6K
1ASQcQvolH/Z2pkClqhFlzjNoBHrpNcG19DDP7wQsmkL1PZems//zjCYkN6CIzgXiC44768gDxgM
WjQIz7fO7Qqc2Y53XYl6HCoByAxAlPhd9gVF70/9VVWqr422fgFXiN7FUifgVWbXFtxLLMVj+aeB
wfaxoYkslQdSM9u3WM9zqz7fL3gWoEzqmlj84X8WaRCIuN0xL56OPXRF9k5P3ctuvhPGrD2AmKOX
mReRzwGxLI7jLTxc6fTJmSLOGUKxCHfV+pjslhTkTHDG61NTjbro4RcigvBIsIGq3HTa6sw5VNMs
OEBNvhTdDdKcRjUJaDjuHvY0IBP7bDm3qRDXCUnrwDZo9vxI8AEnIqYsA4JVJYofYUD80DKREtWh
GIv0ZrJ4rzMWViFuPh4BlNBL6lpSGpB4SyZyfi3H8K1ED4N75CHAtSkgtYW+DO4nnpNKFh+JWgGB
huOE/zuIFB9pkLeqZ4oH8S/5OWnJqHIjvosHa3lz5cNVz18F3UNR0VPPmkssgvLnsYRSkMCQeqfl
xddF0YfyF/bAO69jKpn3RFfK9KYcpAkw89p1/DOfFt9Y07OlNjwIR0v5OZGHsrz+TH2X6TwSD2G7
OL7uEm5rHFYLFZm/wLFtaqMcV6e3uy0MZ4Qyi9CcqURh3yuh+n8eU5cZwNFrSzyzYZdxs791kno2
uP1hV7lD011gAt1euF/pfdshLO2O3hsbVdrHtpvhcf3v2V7xM7qOwxnDipNQjJNFqIjQjV/yKar1
7tnn0wmEg4bd2RwI6TkMZ7UZbaTrkSaJC8wqOOJ3a1KOaoqIm1fEd/XWvY0nMzIWwpoR5f88MPoe
T/xsfjXxvt8/qR2oUwsKOXxBR65bqrLTSqKGID0j/5K7Lx7xeOvIILGS5KD+7v1yseKvVJo+o1BD
QqOp3tBcUdGffjvfDORhiqUGAJszvut71Iq+scHL2DZL9lSy+7t6o6i20j+Io4+cJ0wUd0VsNWMk
orjZxphnHh/9jqjnc2deOd81H6wKXrVEWa8dP/UU1rGGaW+vIqzd5b12NCBHL353Kkli81daVRY+
g1IQnoQPP76YryH4uodDmUxwo3RS+i5ba3SAYOCGBGoE3XxVm5Aut9GjR+kcyC7Wwuk4tQWH73QF
R1cto6+57l9kUWJ77hhMU6tMGveaiINwDRvNcIOccC+Kl4577sEDyKITjPr6mw7gfEBd5WZUqtcF
9P+Vfz6AFu7mY4Q0G6pzInODcQMNGhQYz226421MgHmLp+Sn+y44CGUsaJMkAs9DFmbhkvTTj0xe
pD4WXkF+5RUgsCRXlDKWvdCWjGrdh/uYbPe/uHKVeA7ow7egGpYEz87t1R9t+1BM828jw5uX6X+3
Arh+xgbzvHgG8otkkHN4kpxAQhLQPLiPs2GjKOKAOKuiK/0qXJZDZHiYA5R8VruSCNnvmp7YOBxD
oApvf0rjXU5CgQ0a+co2CsQkwlUDj6j6z/YsMMoMtkXy/6Ul7UPcYpI7ls4prXFY3Yw5F6HYYGUS
7tzoL+tehkcyPMX9ItadORM9Xv9hP0QBWGkP5n6XIR2hmDlKkhAxnzZZUjJoUlQT1DaJ6t09p7DB
5/8nS0+vQzc4zGZ4IJkMk8w9/Bg43YS/gBKxYHjGvLXO6ZbOtZz3rJDDK2ryR/yOlM6eUvQY5B+o
z29cOT0XySjdBnP5Twpcsjkt1iIkOuX6RPo+5L3rUmOmIi8w7K5l6UywyD+CbF50RzQsPkz8EUoI
LEq1qXl+NwZhwu++YtQTTr79KPusO42EXykd30Qo6+dFCFD0wbsXaJh/o0k9pAgypN4In5JZ8Bd6
807wG39OZhzE3JCqeTWUbEklF0aMfmVP+sm8mFnuYVW7BPy68e9RQn2X6BwrWXmOFdBoRbuth2Nc
dqD7ait4VVZgbU1pcpIp17pv67cYA2bEzjIIE9LZDXT8HNnL7F1GS05eQWuHK9haOJ7D9y3fV9pN
uPShtwnkCpPhqNOdirOKdqBt1X2/LrYXL6A/I75TyJzhUIwdxF4W9dsQ9yFKe6Fvb875esu10sQm
iBCuLrzcoxA/b3YtaxNXPCOHPZhSgUoM2ho78ZPuvAFI7+qDnI4ZAQtVEYBQWF1SqPn6kULNXJ7x
OF3RS1PgLCX9NHQR/3qmZITqK5zLYtXi+PCIQLD9VBCYLyq7ZFKAJZ3PU3Y2FuXE5sv5YwZBDLyv
1KlkwHBHUJpy2F6cCk7XL1NtArb9vpJ7e+TVUgaM+7qlP4MCJYXEFtSQdC6tEDxDHcAoOCXQQTmE
0gwnQlfuAsrwYf/m4hhocFi0QNwSLeWRbUcnyWpscHGPl69QFgAQQAnAeo4SMlo/Qvn/k8S7T7V/
gJqvOWBL+Jd5lnVBait0Q4vgahJs3lFSSc0epHF/Yi0xyAluN3eP7JZGqWa2JN2TX5WMAjsI0Kez
vVAx8cZ26q+9iIc9ZyZJKkaG2e6J6MNr3bm91lh96h5IINm8VVM0uh1SJKqjaEO3cVgebUqrVBg4
vlV1id3THsunuGLi6hkueejTwnjp+MVSoPuWfYgM7wzIzJa1WLOo7SGMXtETjX4uDkP4K5ExX8PK
Tis8rAN4LEs1OO5HbxzoXhGN/KaW4laHQ5gHHiEZOHlLtW1DvFBfMN4tjvjkmLUz2VczOAkQu2Qz
O93HfqGGnQYNOogwGxzIiKZsgUBAF93CvcVHyr5iDAeCnMe+KuRa3cBropqrD9SPz/lkpLpvYWUz
Cy2OgyGTKeHMJVeWtVx6Gm80t8TdTOIiYdaUHmuuHf0i44B0eOVehl8Q9E+fLhexdqKmMEh2jPeN
PxHvv9Vnxkew5eZa6ybrLToTQJXGhdvul7CZsNRSqXgAAp0ZjBSmkyrEeS/kG6hJptjgU9HQs0ab
qhMaBNAFTmoIMOyG0UVgTi8eP8QwbhhrqsK/m2bvkS+1CVVX5BSlj8CJ1W58tNNx7SSQg7hge4Tc
Kcgf0qN4i5vpiTeVv4l0BAfZjyrDeSbWIl0loTcTgG6O1N0ciAOVL1QVNWXZZZvWH19wllGGMPkO
rljvIOgBSj32FyLkxBrFdOH7gTbkHt7gI1h1j2O2S0G6V6JoL8HnanL4Dd/SgPBMLPC5dzTZb8Fu
Yj/u6qNV+CC4sP0WMr1kosI7gTsseXmMuYo5BZb7pi8X+RleFL8zNMvxhSO5uQTp+/Z03ZyCyNJX
DF0k6PKWuIrew7uepcXTyKVD7KmFmvHbErecObPRLyYnx1Wb7uq1kVUOXi0cb1Vac6ESNp4q4Ej7
VPLSaJC2yvLFxi+SwXThJvS5Xzx1KSmRbGtmDRh1iCfkPLeRVCaEOlvGQ7Pznj/iPTL26GXC9/NS
x23VGDE3U/92pw3NlFRGUxIOP3krm+ZLUATFIKO7Zck0277won0ozUp6ZoFJ4TbwojjEvY+Zh6fI
ePpAcpu1LF+SVuPYwA9VLsYeuS+Clp75SBB4q3d4mxKmkWiHQcqtZRsxbcmBz3DRr5wo2ZMhY9Zz
B60LYCY9xVSiKPaCe36jlUTlq7dBqEjiq0jsS6XbUJdcT3gR5NqJCe0k/ZOAi7c9XXETvfIGgf/t
JkeolMV3rO7ohW60yIsZR+UpBvjv4S2kEYy3RaIq4A53D394N+lWFJHh31/Qwe+8bqWuzoas/AP6
mEcboF93H+1Mp79LgENkLhuaG/oPuw2y5m5T9tm09XfwVcoEZFPq6Yb73IlfDnGDu2UW6X3lZke7
wyyKLjUJ/5zf5DmQUg+WdVrZSXyekMOdQWEhT81/5y4Lv3MQifEyVS9UyMXifSsdsbSNqmirVb6K
oo/MXGgw5igSJ/8WfMDySExbz5rxv2vlnGDnctk8pbdUcLdyi/t8A1rvpJXIWFNrLHEYMTI+wmwJ
4MSxDVmnZCaPqyavBNQuRMPfHTXvWhoGJj0TSDYRIDIQ0HtieFEVooLO19K2+FexZ1AoWcQ+XwQ9
ik2Eray70fkiAiQuK4FFGmJToC3VIbDW9CGvMbwRVJMfKg8HThGxXLxUYkakq2/y7OF0nlQrE28F
CGuWmSBRUGQfnFT8/Rfw4iVLSu05qrIHVCedr1bI1IUX+JSsXeAlO0RC0+qinTKM1a9+WEiuJuJL
CBt+3YtJHQFJS/4rzhqb2jZp3VC55zWcYs34a4WPAxfXd2AjG+3lM2UUhoQ0FCgbnDjfSfu6pm6s
VYc4THYlWSytG7NFFHdx2OVmXmqFffLpbmW8i5EzvN17c3tVOxE1413XGmHAZ3SEx4hwOz5QeunD
MTrxS+80zgDVkrsVjaN97gjY1QvE09W9BwuB4wO4QEuLu7tiUgTw5PMqcR5hb07jwT42WiLXCm+L
hUvgrsbFqnzh+8rk6tury6DSVFuqI5atXyEUMNsyPmcEnPbb3ctz8WfzQBILKf+IVFoM9L88uAta
03a/w4/PmheYOd7pcLGNHXPC8e61f9zN8yFv7kbUDZrGiMDmCywUQgii4WTs9UP/dRqDR+0bxkxL
IKna90JJarHvnb/EpQjPk6FOIVG1TSYj3qUFDJWhvPZfO21yfynCUHHxAf9bQnc2dhGWc7mrWHmI
Dk4cIVXTWP2bPylmX//pBBxgK/oGizFqSDGDFA/o0nFDrGKGcotJC0QypiFrMyhE+l9wY/sjSgQ8
rHfw8UaQ2DSw5XJGLu9XJ2yEoT8k/rQamHtS6URaR9XmnrobRvXFMnjj7YU7WQFYFJi+ygLDhPxZ
3eqpRmnKVbIBkzLU/zhmQqKaHPuCMpuiSaQOrllAKrMDraQnGmrHQWGGsW2FHcbVgIQkXkxffrrD
y9UaU5qh30HSqE3GLRxQ/DCU753yvvLc0QPkAstI8HdSDFEaTZ9h/Oa6QF/HdvyW1TxVe7VUlp7Z
VyZAnaelIXunbOsz1+PH1+WJAwRYOIRDBuROpO4xhQ1UXfQbiuzUkzPfphwtXjluLvwwvKPPx6j/
mmlvoe4ITFFq1it5n/hpdiHsy9eiDiJW1w/WSKdJEBx279PbkgUcKH+qOJzd3Fy3P3vnDJPLy9VB
oB0HMm92II5QQ+YcHAoZYiDpClO1lPpnk5E+92vCrNE9CeRFhmTgrTYHt76FdUhDMjoRPf1iK7bY
P7UEyYa4gyG/jfIoLG1MYLsWlOXSmJDPfndqQyr6NiKU/7REW233yrivxiQ1tbiBA9s1EQBj6S9l
EmBelVkGxbSSsBV1iSBhJ56HOUT3aEnlj6faQvCtaf84/sfr4LR+jpFJ5ATHxAxeQuJ+l2d30Xyd
3+1avVhuD3pBfczaBO5hOC2zwowJeN8edEBXXGQ0ZNvJQp+PRIsjSXQ82vQQptAW8GNXCTnsLth6
x7uPxdt7moXOrIkAmnSQ9KJMLdvZMhJkc45Vh6gsXjZV2S8sNglHOpgUZjDExbww0HF2DOEKYU/m
dZ7Adas18H4/o1O0cxLBBtZy09VSgFVJSnIYKugniN2JAzxHwPGgw86EBGguQxFi9i5+j6LsmoYm
0qsJ90yiDoHhCTlqRMCpmoaHboUJidmXHJtpRs1Pr60VCCxDN4yShORJOzb+OPMvkYpg+JqPc8Yl
vU7KYz7a8PcWxhxd5TmszP0vVcSTXmsjqbSwNYkAbZUdKPeLsP8+syQI5dmTWKrwy+Qshfa63mYK
1o77Ks9CnC71xO//zYlT55g6C/MKUlco/AFrI8qPyssmrecdYWOyFOKDpEcPFxf8f9joIZl/qULl
9KgMTW1GYr9d6eeLyhj6EsiRAUTktHIexvKTZ5FXu49FgFBnoNDgd4hJV6oUq4Syqm2+aCsOdbqf
hJyRbwTxWLXTstYNepqnnhGy+a4xSZ/+QssyRyVvRqcNF+C8MUzq2jttunGZkGyq0Tk2LnwKfhem
sYuWLt4WoQ8mhzVcm21ANaX6pXn8iESTNEVAsK3iI1GQ92aKIbxrLexewoCua513AIoKWs4fJjuf
eZFyRLakVmrsARoJM8zjqG5Q/Ryef+HCD6KjP+a9PKfo0wHW8ert8TJYofjmNj7xTQHiiiT4vhOa
2lL9YEEFsAdGUlxsI7sQh1bpnNqMVml7RZYk1zaiV302jMcRJubBgTmAVMvhlkBbhHQn431lhfrH
Jm97Yto4RhIInI4MLz1FHJtvBIs0fG8BRxGGdjd5Jh5CV1WNz3ceFpGdi5EpoqWmg00xxytOMRrL
cLQ5D5BpqDpaucEr0cIA7/nDAfcH27VYXJS9EPgxRnMdKjHzEv1AGJO2NZP7hyY9AOA/4EhqDJzl
hFmYVvTTYxLMHAxEW6ye5VgQ8pb8MtyAwOPlcpsv++V8AqVF1Blcsj1foU0m/LjHvz8UoFEuz0Mc
/L33stjyc1nDPFg7VkZYPvOofthWmYNMB7e2CwoZl/F/I5ItDI2wltenqO9tCwuzv/nJnjYPVqGa
EkFcLAP4CAu4p20oLaWMOmCyDibZmwEhLKihrDe2WKy0MP/UW3/idVac+VR13UW1w9isti8hAvDE
2qFSPE1vgFlqNmbQYLDq8Ogwa6DnNp92kR3kBsbg6tQIhwgO3UydRPSOLaTi0vsapH6zhmfYlRWX
nSW3vkfF0zjM0u/Qat18VHSwoVGrQRASqXHnkckf0O02/ei1YrLaI1qnfTsE44G8A7e2ZMQP8MGw
YdNp/zPRDAL41/UUcV+g+z62TuddOlY/nkzuAgZDFBltu9kAgnuwEoFEubPLUAP7Kb8KN93Chf4E
zSrZyDx6GMOgHuYeOdpW071nRlkKXM3jzRg75CM/F5SGIniTYv+cNBKKGn256gR2X3L38R9tEI5N
QugMK7lQDiT36phkX5Ah5hDogt7e21TrpKf+KANKrOBUipVDtWNhqlcybfBGOrHSpRe4BXuSDd/p
h+8GyuiDZktdiUjZjScTIQdoafDb8qZ0qk9KC/Tk/3FmRrgHfl9SAEcMzjEY56L0qYrp/UUgzk4X
+N0q5yKwJX2QdJ3XKeb1J2SYB/lR3ayYzXgODm+eX8LDFEfNbt6VSWiTUghR0OpzEUkhVYPiHU24
dgVto3nz4MU/lgZMuRAygiMZxGYoqjaSxKcOJI1m/TD37aORMJG7uQoy5CSoqC6EPfSi9vddWa1p
wxt9PmVB55XhtmjDaayuROVNCjMCvK6FdTdOmP0YML3aVappTVO5kpGyIoTHLXOWgrol+zfRDui/
SCob2ImFvDSh3RxsnD/i0wDcH/s1m4dKGoYgGk/nGBY4kfXpjqE7QnooshNwiWgoSbvxhH45miH3
pF6fLYU4KjFQUOA1KPS7I3faphykGvAn+k/EPTAWdAZfaFQVJHKoXyFsz5dz/pZLt4qBR320Smiy
1lDfJkE96ps9Ps+1niTYWEhTEFoXPeFKXv5Dq00CKP6QQZIj1lz49FgsIutDtYmvsCJuH0lbVZ3J
tp+2Qb94u6qd3YDF/ghN5ABi4/9a+EQU3elgg2bMylfxPXLKUaMTEdqn4VKNRBvOqENqGFWtr2br
RMsN9Wz8UTMHaZuHZChebPG9Ti1h4y8vREMSs+7hS9QLh9PXtl+8/v7TIQAKNakt17gdjARL5zMw
d9GLQRhhpqaHDygu2SDH7QUYDWIOxCqR3lNKXZw33vQXo3DrVU8RkE0ol62zn/wudQbKdxp2tszR
+JIS71X6o4LTC0hDmAhoPX0hwp+eLWIIXnaMaUGmaRAizTM+WAYCZXUA6rNp/9rq1ZQKxMriSEqj
sFxF7zEYDVLPSmDDiPVRe4tTOyGYkNJXSd2JgOS5Rw9DYPY4Aunz53DMpmh+Lz8FT0r3wNhipl6o
/bYPOIEKu+1aaUHEptnyyxh4ha7LjDiLlWrJoNeUbD2yFnMuxP2BeTru6w6FVeUtdkCdohinP8Vh
u1O2nLKoNTnYCpGkyD+h8j25wf2Jisc1akfSWiOt91eCQcR5VqR0WVAzZS954CGHT61Qb1As+qs2
Wqpi9cAVaJ437dA/NVE28CmISRnHoqxvZ1/LOnNH4QJItqlH35PCsuvD74Q12AWDq11cmOUOdQYI
j1gcVxCQwc9i+ieELkOs876AGO4CvkaripeDumz9maEa0JwSzBdsfs2+8lvYs6wC7CvooZRbDGJY
yoLH3QTvx7buJrrLgFyYyVnWkmQmXau7DMHD1gxbSTVHT/qrraaUlsXOPWSiCjP6YKbA7a/GeAUx
2zIWLbmYD4thjOXk0s2Mwu8HrTkROdaw0Rg0XKZ+H5saJn2oILGYLac/Od4a+8dbuIKxQITQrg/5
0RZoy28imjbtuVgU1lgoTlQWE9N+0mTo6h3ISKG3qbsXGqvwnsM4j68UgpNTj5JzUqLq96n3iYvQ
zuOG8h+L/WpmHi+ISJvPrK1ODACQd1yc5+Rfo1kL0ZJ28LtE317AUVDNp8p7B0lI/r4SI+PcrsRo
6gY6+2P1oHVZbiSqxwWCyRtGWT3e27VH3iWeiuE5zvb7MAPbUnhDcNtkvh8kw/OWrRW/RVxk4KsB
TYfTDr7mb+0RopLhZx0mVQ9dGFltTjWhhcZU5cyeX5NHSy7cPxuuCK/8ZkUEzZISOr1H4nAUq5SM
YzOFUAU0NeK2nG54JlgYlNrEPrFEm+UMCPGpIz5BGkUwVwYF/wuYS9cU0e1/G86Ipv1dhGLURljB
IHsQp1zISqIAZiwUiOaW0p+a6X0AV1rgfkef7juZRvXXMEslQOlY3z9aw17MjIaLus3i6o8aiP3Q
NoL7pAqG4ru/DVQ3loi5lJdNZH+jaeq6v5e0QgAjtT0zkBj18PZ/15WScNupBpInrphO1opOkUEW
+CV+gz3ToX/uwpzlQyD6DjeRxKWqLSLRhTIek0QngHSJllKRrvt3Wvi8tkXM17iOhZ5lIDroIULZ
eNohWRNIhwdWcwqY7MXRuGm8lVecW0W6bN5UJIkx7bj/tfbf1ZgrYDdZobQFxjT8pUB4pz6G7S41
yb46lRqxFT7RU0W3A1g18b7iQZgC4JPm7cbawYo26vilKQ7BXfJN/eA7s0t0z2zcWEhhrN012X7S
FYw75gjTcAeXgvoN8azGIqt3qzHhJs8eQ9DX/auDZdxLKci7NpGJjtEtt7rMynHpnb+huziW6KX6
PIU5qv1FWYguAJwjwuSKuIjHst/zp9wcKrDJ/yxEOd7uefK9yh81Hr032c7EernXCwARDmYkcMfo
GY2VFWYX38zGKDs0XAdeLoRJweFTA2Dg6kzU/bfIKPXfOXrQQx0z2x1IGCsc5ZDwr/Jlc5LObR/y
/5ZJFDfDznscTcxvn0rLmYa05+u/G7c2GJMzHCAEZmaIaDo3qIiie1JLHHPHIk+MRfQ35GIvBNps
XVVKlHb7mXKYBDJPkrNGPbBoGtpTcwF/T20hWXLz2lXfYoYg2VVAcBywFuznyuHACvPYbn0IA5lz
q/gQoWuWsSUHtx9Om1eNqMfQ+B0+kuqIp/Imfywtd6rBPtXF/JBcNAAm7/wyMqx14Xkal+S2YAyg
6gm19eUcUX0k7erPT8DNc9rtgoC7wo9fLKu/0voUBKmkKKjDxzXdZ5a/jeePq4Khvuq+hDMThpT7
GLzyZFgXOmgxhdOcCdelCZNYsJSWAyrip2MHaVVfWHgC8TMJ1fZPa0rfZhqqwK7QQyNuR/UruKu2
G3ca6puD1AwMjSWqyl9xtyzcuOIqm+LyhzuFseUje2FtHuosFHFgyulZT5JNvbnquAukjWOa1qtM
dd03sm0T/DuwQc+0dkDxZK3s9Ie/bc83rbIfImvfvhhN0W0TW1UyYqaqCR8m7tHmSfeQ8iwHoPbf
833dNqkyd6gDRR1qnt+mMQu/v71M+6H7coJRYMLtR0CQVAFadQ8+Bp9kjnkHHIWXBFaxuSQ9DQZq
nQX60zNP93VPz2arCxMT5oO/3q3Zep/ZqPGkOkXVVkCvDiZOUJ3PhU4Pj497mLnf1t7HodcHhgxa
a1gcLS/qHQwqghpinqaRgWz87m5pOo7S5TrP0h2SAbWeWsnnde3Wnv9b/HeBmFTjFJOAzsWispkj
I34nCviuBQPCLO8q9GhH/t3/pVT/3eizdyqoBAGU3QELWA1kAqChMw+rcx9jrvTwj7+FOsdlNOKt
nzycvH9HM4JdlNJVXJBMa1pzMmBrgN9xQJGoMzty8bXrK0uqXDsLwplM3dryjjUAZTGWrrrCuQKA
G1dyAXNRKhrXvFOVG1KuRGaFwEZXYZiWOEb+exGLCW4w4ufvCww+D51WZAJ+/0lgNBFG484TG0V8
GzWvzgyx3iyGTiwN9WNjUjLG97wpuB5ESLgRpt3KLodNQr+k/S4MemLfc3wbTfpHQVmJDSFUwKtz
PrE66PbcQ2QkpVTfICPXnky9ksUugdfvuavf3fw5S9u3lrAlGTC6w9a4gRsxzmWi9scidgmUXpe3
RKXIad36UbWMusH71yu2i0vgHR3OeoaDHbNu+oqNu9HG66hmpsg+K1eAILup3Uw+DTwTqKz2lvD9
CAlfFHi3Z5GjSinYszEuwtXAU/W8TQksqcrvOn2ufvh+XajnAeQMB7NpjCpnjwYS/Jd/qekHW/QA
oRD2ns2kzmWhUEH8SG3vvR1jcPJt0Mytu5IAg2BGbnpLZzhy2zh8R70Q8OlcqeQjjyQRk2CmYlHW
bzIU2bisitdpdzvzDmtQBe9BGhjge5MebfphuWx/CLKJiBvYCWYaSYA7Vtnb6a902Gbra9ZkJZ7i
A98Y7eJg3hhg0s25FtSoi20tP9Tauo1kdYQ4uXNiNUNPOoT2ZuqK1btT4+pcJIW1qQjjksDZi71s
9ow6y1DoBYT8ja2VpNcda4dUaFvlmLH9jBuXDT5Rhph+J8gM47++6TY/VU0KVoY8cdLqfWgKNb4g
DTFJOabsJn82i7euglehdRmNPLYL2tUQRnv9VZuAfNlU12JER809beylPsALSM8lBaT1tcQIndFw
5V4+yB5lJ67t0E+XS3GiLyHammtZIAB+dlhjENFY95iKp4kih/GRf7tBzFIkvJXwci7Dm7Q9YF+H
Kjgrr5rDnWUYCfknQIhlxmbmpUT5id7A6lY9WuV7e7Ukq4s1/xaizmrfKGGEdIMy5duRQUqaeD1z
+5uohHAqzOC4YJ/pWFg1FXmNf61TgvPNamnWfyJB9aikbsBUVI8c9iTbyYYBTQtfQ/pIkSqzRxT5
+2gPWZwf1k6G8TSxE29V2L+PoCBnGv3ikPtUohhJ+zW9JkFRCY1sSuh2GWpfFSBuJfQHg9kV0Obt
+qXHdBr4VP325xQrIndiYLTWQKyMkmrBPEnnlQvauIlMO/ulN1G6qbrnGAV+Vb9PvRBxBB1UgvRO
3ZIguXA0mC46equX9MnQAsVKxagl+Hc1FIIE7bzhdmkfp20a6YZky++qPkCQIvPc+zMmvXoLClhG
7nucKEFWf3AM1Y9FoEouDhI4tAArhKE1EekIRgKseQZSnw+hryqdHTlQ54YL3mCPBJ85MuQ826me
8Eu3DnrMC0laR/dH8V+3b15lgKH2RwwAwL2FcD/NgBlhgf58Ijpff5OjelvqkqG0M7AjHdZZIFxy
3ieU2LBJQ/DurcHP5gMUF6jYnFRm7rHURUUhIRV3YFYdahNpwM8MZTZUyJMzZhqh9GNVCmFrS6K8
1BA5PTXzaYLtwm2fotzrojsAcZ51CE8XvykCbMATmpQmxFRUUg2itVVDqseuZMOvb7sJ1803s+8d
emRwjBXRftRXdDN5VscaV91Hdst0H7m9ltZNOWguScmQpjTKKG36Ge3v1++pf27+Cqrdh3Z5oSUz
Q2ud27FjnQ7nc2jMGNX+h4G9G7Tskdf7uTPM3qFtZBYUYnpqC+DwLTQtcB4gcgRrPvfUkgPT0xGM
V+GGiN4poUe2UUT5sX7JHiyz4litluU6jN0Gy3efkMYTF9ee+XlL/nmR0KsHmjN1EavjkVfNyZyn
VTZSeC6FRvHPVyW2osawQMeASxvsuGgadtVSFGOBkVuRlV8ADYfk3JbijGHGcKhbM3L+1lfDSetr
bbKFxxfssem78JkTVgRFBm9WcykerpgS1iSsM2RzXaejdNXMQCMyBKC2LyVggLZgZBNMT71roxgP
XkMmfwNcA5PJc08LW+Ik/HP3bg1EFdmLdolQjTbCuAAqOLNkVLKFn4VXV4FPcKZQejRI4qC7qGjq
i3mbElgXKmbD+4vIzoCmZWysR594p2JXNi8I8AM9UGynszftVSYOdzEHSnmXveNSO/WU/hnhl4zh
l9dDWTQTUUquDPeLc6ZqSBuVoWspYh3ECnOtoUB3FmgBfM8Qv7+OuSfuqwNMWvwj9cUIQKBLnhjg
O1WKqmtcs1qkcJr8B9f8Q+ifG4CMgtl69er42RUTrmu+i8gWxYg9cNkKSMBqWtRqW0169pYyNMV5
/aowJAwITd9CrY8lDUmvyTyIrp/+QBroC6dRxFFL36js5Z3KKJgZnwEVj+juG/ef1sOHRNPu+5K/
ctYkNJ/k62P60Mply6ZFjvQBfwOJJBnkhp2g8kIJ9pG0W/ATNsrRDqzqPqZN3p7HZQWgCwx514YB
hEQ+G7EqfhSMvsC1pn9kfjiCQHa7nLgGFcGp8K2yDIxRTCODW6wEIuyqHiF21I4TPRtWxAF3czRB
IQP6BGoPJLo8Xy/zgHMIl9Sf7FQD69G6b3hx6+BfyLrlXkCq/xAJDZA2A622wZSaLCFUQ510psKO
X7IzKzJ4m614V0q5K5o93MXBodKXVVyw+psz4QD7WXIfP9DNzs/v6ori8bAa0Ymniccf/A3hmYy/
E3lwlLZgnWTheIdVA0uY+MFDvvTU6eYuyp8apEOgIB4Ao1BhCugg/gEMkMBJKmBE/nRKhUBAHawM
6sbjVwUekYotr0KQOQ+Yodi7b14aNus7DECaJuCvnT1lX56EtKu70QjEELkUkPt6041zE7W0XPFU
sOd5mSP1YmFPbmQSrB7l7NnFedwSdls8chtm5omknTVtJdEwyIKGlMY+XWtuQGJwEhxM5/QWV+yk
IvE+VqIJtiIO3ZuwWXY9BTaQJF/sFTC0AiJhCuI6SRbepejkV4l76EJ43TyPVcBR9hs4e1epb4K5
wYDtZSNtxKj+cJrRglAUAkMJ4Nf7OxhV4MULZYtkVlffIXV5oINlKIYYQrldBcwyl4cBqJfc733l
ZXkxKBdot8C6UNCCm54dcrPDQb3gUPJdv1PdEQLajpvI2ynE+nML/j7VD4oJJfCzbIjeqnyS4sqK
dlXxKkEkAgJBMle7RUjKd6+8uPpilDoeYuFCJjgmaVuKjQjA57SNXFwzisYW9mWIk1V3DPBAdN07
6cgJ2OpRZwhCtYKz+eE8xyyNcu/aiVMhILHko4BeOwXF0s/R84G8mAdqKkbJW9HhfaMrlrlVqdzz
v0qaQfXG5seoQw03QtU9BDwVHqsZ7EqPOIHIrHtidQfnV+prkGi4KWcz6eHdAI6HNIfL4la6do5F
d9LEIDJWTeTKdbp1nIXLx43vPTut7NqVYFcyBQoKlfRRr/oHFhRRnEZosG0PlQ63jFxFIITrvNAH
MhdH3niyRvK+tPt9MJ17qibsP1U4jgycZMVZkCikcZGYHoyEo5ywBuLZNTziI7XzrjB64sZWUwCh
lcjA/Z/HOPfsSAUjFkKi6dBUIuF48rJCBKQaAVKEW6ZFljPmF5d35yiZ+srUXSd7iNqkZFM6ExSz
77AeK+JZsj61tP/2fQP4vm/JC4c/G24FDSfM2fZ2Z9jaRvNvnd/IyFpQ8vO/1kiHt8VlkhuX/fhj
h50FR1OAFgv8qzl5HWwRu9iAyZz7LRfDzBWzA3gny+ZS+gLXBu/ev5nolyFo2YNdKlmAM39wIDPM
lxnFpPaidxwtxaz3H00dnvrGG+3BE1QdQOKXWGz6eOCHVJrx2aCBoVl03RLiHCCtiGd4pOqEi/q4
rwK/QQlAogMbxQ7r2BIv122iVOTpK7l7EqHnAL9cJNlIB5b39AahCtZIR88JrJVy9uTam4u8wcd4
A+7KxYGpEBXQzo3SbNsIOzVgJToOKmLtcl2wRjENf08Hld710+VfsAgv5+q9GDXJjhzI9E4/0hAD
NjlvE/eC60c3/fA2id6svg2552UAmkyxoukUv9oRFmD4Us2XtCOk4PqPfebDG+c3Z42UxQuPacQ3
xYFLzNQSY3qdJBtFVhipXmEVVzvagVvA7hm4U7bCaEG4/4o53/OvrGpz5XY0DGcS/KscsCE0uv6q
5DanyXykxXouyU2fJdulthpYU32FcIlI+ZfmFU0TlyfbSITpmwDOqczuyz0L3Yg55votWCGKYoB+
VjvMDkzjqh9lEYAVPKIgfA1dQPNEdDaakF4XHVl4ldd3L2q9+P/WKMC0YsvmIZlizof3wUuaL90q
MB3ItsjP3KiyNWxMwhu8nJmrhH1LdT2Rl60QSKKJCAA9WfyMZAkKPyDFgVnK/a3AgiaVixPENPuX
wrDssz7Wq2turPJATqNvpcXeVPI9Z2aTw5hAmKG20FcPTddYwbP22p0dRXnEVxGspNjnAEXGmbK7
hWgo0NBXOxxO+MNLAnqaFxJVo/mECe371AvGKHtRutUJhEC2nhXDkF8eXCptcRVE8COVJn2KZCMp
OMLoiya71/XNShP35PKDozl+BkGwY2R67gGaEIg6g17FWfIofAFCw74rN6HLt4bRU1uFZxKdfjCF
SJ6BP3O856Yj/VGsOgXUxn5HfgJ+1E8rG7JAX3VKLjlbWeRXikCN1naXOIqXLAxFWs02nFipjkyZ
Xd+4+G09ojMkszhfFjAZmsPiV4nmhwJ1gTvOcQT9p2QmZm72AIwc5BYxEQBcdNou/3vm9WQ9tgmM
3L+vrV7KxtmFu6RkqHVzNPvS2lYiA6SK8xfNm/S4AN8o6muvFQRlwoyyBJ/K231F314Z773c7KqP
ud233Hzbumfyih6bLwCRz1J4gvlx1W2mhHH+RYWYmWsMDlMP4xLE3thYwQus+5wwgxcxV+3GB445
SCdPVLCg0ZyXArxS6fBspoQZ0dra+zLAK9tYz67ywR7tHdAgK+AGG7xu3JPGzHf7nS9Xe9jP17+E
mvsB9SJp4r2NWSgAINMZPbOL6EeJvZMTpPFvna/gnHa01Qz72KVB7JpxvkgDXrYUbZdCVeqAtbkW
+cP7aYRH5jWe+Mny6aKHUjvgoadkl1btgHZG+HD7owx+/oVwZY1FOvZs8Tq3/cnMfV668UzRRExm
/gds/0liw6qkZADm4qABxRW02VhS5f/Q8MEJiLsDexnnuj72c0623BxH9TwPnAyxm8oXQDwdUJaa
HUtn322DlF1ujIFw/42ZQ8OIKIwXihPXDNJZxzoDezqLTHbzb/smAyU48tHvhjv9NegQG5GsaYTb
dfub6lVB0n2EY4kRCifz
`protect end_protected
