`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fbDaBFHIKh52nacy9jMzYCMG1Qperci1BNhS3a905yYf8AeecKbmEQtlgupMzzq2Jx4PoYceu5dv
l8wFyM1beA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Utdt03S3Lz7i7p6dw60Xpdtn/qfD30vK9yxGkNw8JA+BhbYYcx2eoy6xX3s4i04F8mu4ZXW2yaRZ
QiRt02sJxlPynHgxFzZFQmLJ7VAzJcFAktOKXhWNwj9wLoAbrMTsjoWkKcK0jFv8BD3HlVd+njar
EYmkdb69Iz7LBFGQbpM=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4PT6F7RUlC6ulkKy8EHrmmm//6hC9n04KErb4TQM3+Jh/QcJmRo2+sfuzcdUkdDM5tVLyoL1zas1
82QYOJGjRNqJG3/ONBtWFb1AfoD+7KRaeqKM0ekCCP8CRxqTvi4BLAj7qKoZYocNy+9GHsu6grZb
IcibNZIQIW4p5GlkwaM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oXpOej2si6vfmCwhxT9L2hA9y+uHvnEYR0CqR0g9lpI35C5OC1domnau9GAI8KKsKod2cMYkrO7N
p7BfJt68O4gx3HP2fnTtvSGQPi4hCU4JENf3ea0gZptV6Uug73DvcxlphHzEsfQvNDytZPzCDl9i
TYJRC3+nNJ17CrUuAjQw5TNZ5CEr0ab9sR5vNiV83iixbHVzhRlMWTba+N49pyQq7xLXTuw7KA6M
WgaNEcIO3uhOCpLBhnmF51V4crqXW3jbuHGHRN41+3s4eLXkbwxVGgIXBKdxNE2911IrZwlBIEVI
fGVkj/T3llHvdFKE2enmfnBtG67VsqyqSxxLDg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p20y5FqSsxVqxQaw6mFQUmXW0btKlvrXp4sdgMO5NU7I0yS2G7wUu4HdQz9aEDl9Vee8yKfezePv
lKk2Xic9pdtgGsPnB+DEqIub2ViadwY4ObLTLleVBZgq2zcbDjSiOGkRKMcizquTL5/BcxMdOLUu
02Bsp3MFcDoxOYy8ciUkJiA5G1i57Yyiw9rCwr2Ta5+Yyi6RtbWM3lm8yQGLM4PubCTG8tkHfClF
WpFYFE54lHbdMNH+GNHfUIWynJ4avx4pyymRgZ/1Csh+uO1sG+rm9LtQ+fJIOKsR4UqptvUtNx5+
dQXdpnubb2XNE13HIgKarr4vtrXwnd05n+buJQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lqz0XM1L5SrgMWZTZt3KjAQO8hxce+rwEG22w1QNMgpWvLZsg6hKjbPLKUTF5//u48F5En6+esxI
KuJ8xEbRiHqjxj2/3FhHbQyfyNDY71VV8lk2FNFJtZH2lFJGOj9F80zlm3kmvhwdLSnrMDCci0t+
sOA1BiYTZJvdy5WvwhrJhOJ8uGLujb5oc2C8InL0jxeZPku4c4GpPs4ClG4Vaqujl1YuTHw9nwgT
2VoUpAezNIeVLFOBUSIkShA4NcbLqfGZPQcX1fNAoKz/yN4NE9vB82uLm5W3b2B2JjJoX2c1QSoK
msqvphRnK2MpZEXP0f4zktg/gfscI47gPQFk4w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22080)
`protect data_block
nyGWB5qqpYafdnMqNNuNaYBWiJoLpzeJV3cR5EAujZEWREaXa7f7X6ay8CELAUdvsqZTqugJYyqF
1znrpJveMvupAwj0txD3xOBtOEJimn6HymSm7mKt0pqaIXQ1PKyKfY/3pfiapUfarNN4u3RJUSOR
6jBTDrGuMM06VP5CrgA1RIYl+LyrfutoiGjf2bnPLebKVn3YalRcBohCuVvSUmDB9waX5nrpyRVG
lE6nLGP6fWIViERAK9VSuUh0VQnITAc4/YdHI9iwUpuUXVt0WaLD3pXUSFaQoz8fLz26NufN2X5L
JV23tVfogUB4GUrv46WFizmNg8Ym9JrFErz167fx/jyDbs5+HDkDYQ0s5A+wge6wsskwzShhNMzk
9X1oddNZxUC6WU59AES/VHlWozplmd4EaryoE6f4BvKj+kTASTfnwKz9Tmg+vLb3NgvCKn1MMWzr
MJBAfPiRinAAdPcAcZ7v+W0zqlTAjajs8sEDHpEvH6EXY0OjC1uMHHb0uiNirCXE3tC+5zfWJH3e
hkiX1DBgqbTzvolcdu5q9k8mTlWhV/+WQS4WS8IM6qMFGjbxc6urQsrkcfubC0QcU2gOtrVyJUQb
6VsVc4P2yNZViO8TV7STKqYgSpVSHDhRrduCZtVGaH0kZOWdtXX/dsAZWiS+0RmvQXu30K8QkITA
SHICV4W1TCG0Q/H4v2RFg1QM9BhP/ga+LKKJtNic0c6AATv0j9EHO2ruvFHT3scc74P7CMFB52MK
4n/qKFxllKuetjeexVppArso0gukKVgCacbmtj5Fp9BZvVvoDBpcPnmiDDiDyOn9W0BgwGSCFpyM
uOQ8V5TKo67ZL0cvPkoaWAVohVYqkahHCSzk8+USreD/kgiNfsXoTj9iK1pWIOGDDNv2/GSTK7N0
eXVeyB3/WXVra/s2xUK2Km6k1+WFQc3NFuqfNqMxj/fZbW1HOh6VMEV6b43dDJ00RTj8jg5TKDl6
aRIzX/h110+ZipIIoY+bjBoAIj1eeiUDTa1wQhut2ED4bTG4G72hONa5UJ8RCAhSnty7ofhrWEtJ
OfdO3UMx2OQEPDFX8hIVbYxESLLaOqHHssZG4bHhKi82OW+sUpBNv+0dpGNhrppgqnAxwGtF+uBl
VAZlESggTg/CYe7Gmy1BEtc7vZZTF0D0BxYkAl7scXBoWVHK9sKNNHM7VC1Ht45xOICl+fyuJmWY
g8Lj5T9WMeQVxdxDIe7Is/L7KZTJTH3GtKqmIRKiWEAZpP4RY/fGlsChO5QYNwTHn+5l7RCeGpcn
qGfQt06oOrhn0aOxbiZ9D3sdfPDjezZqgpMfc9j3lFGCUpouVxOIAQH2K+eRo5QUQ0ex+dLFR7K8
PmeFsDVp4wPc9xZs5miLwnTIFTNc9CChFmz6RsSErKU4Ft4B9XScbBsq1xIv89CRsUwYmq23Ny4c
NZRq9Fg2gsXthCdV+h94YHvUuMdPFwsvMOK1WgA0SoaqLXaJzZyNigoLnEEumXUQaPkSm36pKuPn
hAQs/n//InJtxxxJm7lypT3JNx/2FpAAKVQy0agAHLzR1ZWkroagjI1yqc0+WNW60PGUilo8HE28
ZPRUaPvZXrVz7shHGcmnq5Yii79O23YMDh4yICkdtYJNQa2YPMcYGjqbu14STcffHUuYNKBcszui
4eiircOOB7mTMrdI+w7IScjPPeV8X/URDYDtLQAbcpB5jdpdsf7KvVIj64DWxIsdqYc2ylaHqfSL
xY8baE5kRqIaiUBLlIMJD2Qw0Yvkl2yYmPsbvFJKjV/Vt7ALDdIT7YHCA6Q6yY2UmU19ItwghZtt
Lp2MEbEObkjqbJfwBZWuVChHI9V2rPlFTNEXazQcAsNcug/u9nki0wepEU60vGnA0YoGvCO+YPPo
XMJSe7zy/b3tD/b8ONGJc2w1drQG35/UCnZbm096Bwf+G0M+VNCHcehhiDnKpQIrrsotkTB8IQzf
KfH2iq6nyd6MECz3VGXhNlx3VLYbRloTD5hx9hE+zZW27X+9tAJlWUOciFG3qqAJlS7NbAgqh3Nl
2EDT95X2ampyY3dPEq+mPrNh3cbYZAHoKk9a+ojfjv5vbnmv0pJbGdntaaxj91Ga26X9n05IlA/4
TPalXYACiUKn+W27sVJMGdIMrsHk4RtH1I/HimgSDOzaxsD57BgetzahDg1qJ2BRT/A2R2qi40mx
JlTgr7O7C/DW8AXL0+BEIKQjz3G7W+LWYw7iZ6GeWRXs0KVh4MP4xAfaRWMwqc3Dp8bWEwnGPgZT
kjrPghDD1YZ6oCDs8TrXM3Rf/xjYmfRk0oj0btK7WaBnm1l9wsIh6t1NxBaxfuA2EBi92HREoNWj
dJIYjjaCU8IysuaMntDm0HRuIt6Ygp4WkG0VWh/d2Z0zmpyPujU2OSDw1/kjqMd8Rt0xqSIl2sqy
jEjnjxxx9BGvG2OBZ5AFNFhR+2cNnwY2zF98TIeGLleL398OHyX66hFUmKEd/VUbVxJb4oLiyJat
iAtWF4btbPgBb1HoeAe77nY3qJY3EHBXtBmeLLkmOWxUQFvlVFUSrxaw4wPidWufsKoaFyvAv9sc
tEfu7F9NCuIR1FfI2Bue9pkNiQ4DWcECOuL38aXW/o1DRw5O4/VDvDRRHwIwCd9q302rJG1eM3Sa
I43bOtS3JLHGJ+vGqC8wGfrBQLmP84GHfhynuWZqHrIgVUVwx62RHTUoPh8Cp9lbWxaMxOhjPCdQ
dvBWuOD/6ZwUd7L6247Zo8bJBdlWfOD7M9bZptl3BKr52TFAEvb0bw+UYO34V7/91jg0e2TmpbXY
OigL49gQzcFpVjqHzZyx0tod91BkGF0NE6sbXAM2DcxiZ0yM3u2Fa9ifr6pHN/ipR4klFuK8ehHD
61c27qfRAf3xGnLnA1yk+z7tQQ3g2ESJWaVNRk/SurEXmrvtQWLKQc/CZl1nPnKdDXQsjGJUJpaz
28nmuw9ZqndCaWitFTGtHtaStzIaQTafLFzpbl5vgRY0EtEQgU121DZ8JmJbXK2pNOnMPjxe/vpi
94WHTfz75Qrxxp1OqS13wA04fAg1jaF5gnCAMie8gUgzK8S5avKEmAOWZsTWthtY2C4AgLPD/KnA
e3kQ9tKb3q1kMfLfNKUNh87u9Tvvj96NQEieIIiHcWtr8gtz6EfCkTCbU3I12YpKWCG5Z328/Xoh
jf69S98C3pF68ZPTF/mv49X6y+92FIn3lN8kI9uX6oTVoIrgeIMbkjqtWzL8Ssyv98TrgsuHuGcH
AUxx+biFAxnPIv9cSvdNU9i0kLU09H5bV6UzOyA2yBDFUPZSWMaszeZHoRPa/XV57wfEkICMGNMV
bqEyd4vEk8TFetm3WG6f1NbUtZiKA02zHxP30qIuFN4pos+sL9JvpavT8I6czr7ZIm6Z61AI6Mhk
U5YdmOffh8u7U0XHmwn7KeUt8gDwbHSu54HQJI1JwmMuxQy4Zn8rA9UZqB3IufrTx4X4tVP38+hr
mQOuzhmMQURInf+QZ7ovMRi3+pLPrJO/ADh8Jqyr8BlY4Yg2spgnMQO1XLGPN2Cx40jN8HbDHdR8
wJrAKkMi1jU6IzvwqNpeyCuibsFGwxr1y10raIGYpzmz8Xmxy9s8l0p78l4MC2BLnHr1nE8koSgb
+t3eVn3o25w/vgLtU5Rv6G3wySISNKRsXyDPRPvVHzPsrEqvD8kqhdc/kPsfj5jPzSZc6/Hj2IXg
YPTfZSRiuGeUB/RPAawVjQapc1oQkO2w5yBtpvDeDY3++qLgttBXBOZgyETKVy/uMezsV9T8x3Pn
dEYBstTcLbHyLouGOzyQJ16HzKiwaSbCUPtlBMJNZdvciGq2ThjxsmFL5x7V1/Q/JU4OA22CefqV
Yr2yXyJ5Nt+PfKNDrXcfXEHGdaF4uKLSLNvCIwQExT4S/Bxkm/wtbhI7TcbfPWfPBqdeuJ5IcfGV
PdjAs0Ef9Rkm4x4ER2l/eqEkxXOW1JjayrvT/IuckxbnJSVle3yBm/fUrY9w7uXzvlVUHbH1CPOn
unI/Hx4EOONUADQQrH7YzTlFbzpk4PoDzai209SGMF5nE7bvpMDikTAfKQW6rbMqrt0Mb6T6QpNL
AEBUfLDdmy3Xm3QpMJq+Xzt6SA1JoUjvFTSvZcWFT9XzvpJ/LJJKe2jWogzUnsQilzeIDx9WYqQT
J/WRwlSfm2MzPkJ8aG61UgybHvae9g3Hlmlb3DfucJSmb34kKd7GSzjCLjQji16FQ8qxtfVO/2i5
JuTPM1CPmQ0wB0zv0E0NuFjCzKfXlmyexoDq3owlWtYfFQV+US1Ji54dMVJHOcAt9WlL2XgcRRrV
Jcimah/ck2RMWtP7hn7pTcT9uvHFoOdhnMJBA4Joe+N7emcG9XdxyCrQadmpRMN+x7/0OuXaAVwc
esKddDRzEehm/nVjhUUtGHDz7cgqgWOQn3sENMkUDLV9LCpjU5GVySJaqbyt6l8tgZzj9od0+dR4
zqxyrsApbRIMN+kcpIvV+WHUQhFARJW3anifQRTjSV/eaqfIrJDaVgwH+LK+wBfuIDq6mvri42HA
LY8jQyIHOQc81iEn5iPOzxCEIN0QeUhUuFzDlp7HdjQrAlN6TdHx1g3GC9phRcN3isVKTuGbHDbY
NKsydKRjdjgtpG/FsUrPay2JGGFlP+KH4K7js1NfFQIwWIqYkijDuqAbQa4pbHx/U5Zd46libWmv
NYXDpb1kHoWFlqpMO7epHPo5dLNT8knk1BT4CiBbwRtQs77WXjh4FNrx2z0eY6tOCdHl/5ZeW0Nf
aFLWDRcdRq/KqsG4qXXKLMGt3EbqF9yEpqW2lYvyBjd3XaXmi8YpO43JAqIBImRvaYCV6jd9FqCZ
Z1iK7QLSJUMCOmQkaduj/W2a7OaA/BZ5qOVeWbJXuj3XpX/xngG2wIfymTCysiVBFYUYSGGsX9nL
zKoZDGqCoQ3WyXeivyw5eJup4NrstnzQnyd6SJSt/tUKAcGfRQXMka34MjcfqfX9B+fhFTHoMiYP
Iyx8EAeRqKvKfyvoG8zylCfannim4JI9fzAZI2GQ9sQ568EdhTC06BzsfCeQZrOgare/82azYhdn
oKZUM6y3P7SBVKrYi+ljnxdFeCnmpXu7j1BxQ7dnZQ1RS+3QH7dV0q7Yy/bNyxwmCL1RHiOdpNhX
GWrB1JxlgvSW4DxkWVALxuJi7BrgI/BAbZvrb5us/AVM9kshkl9fO1Uw7bAuXK/h0n/2fSCY7kze
c5MmuuEIze2/ASfLOwIGtSGSFmzKoefMYl7S7m8Zz0IRFgfYIRHqboYUy6lq8sz5IzQ/VlWPKLqa
l7NtWecSukRAjr7pFU+ELuhupw0OBMtiIeyqUC8tLYdWysoai9MwM+BEjuPrkypT6Ztdg09WiruU
qUlSz/jBWM8JcDoq7K2ifdDat3mo27xsZr+F225tj/udOPTOOnM2uuBP1+yG+jqw4ojT17cZzidg
ihluLCy0n8DB6XeqJdw+56z6vWoxYSKMkEtw1+E1ooXwPzwFB7C+CHSMIZTE2F2rCWtZnTlcv4Ii
9l1TxrOXI+R8L1CxlLAQej0/Jfl4SPIaI3UaNECuI5iLuoEGMYKiFWcsRS73qobhwtsG4w7Ma6Pu
RP5ppRdUFG5bEKFhzQzSYWha9EyGQInusJRXnl9NpjSyTLc8bynWbIUyuRa8E/T61o2BaCJUKfQv
6xyRMajEG1Ky2y8pu3LHlTIJD9ygiYXlbUdXFgDvJ53OTLKBx7g5yppKK5sxd0tlmaGBzhOgXgoL
Ic8baytqsXHMvWnBqiJlwPvuup85+6i9tKa7grvRh8HPo8+hdxlmO9/6SliGqlsu9967bbYzYHDW
Yw78s+hjdZSG4MAYVsjtZBxRMTkWVvTjmTYaJnKoCptTOOfiEQycOPhuwKDZ9p5vU4kqqwrzvf59
WSmral8bPKQEjIsnotsYDxZgY+H+XU0ovEuy+eBewP1diyFShHZiSuLkuwkmLN26Qdgj7fp9e7dA
6CKok/VF50vpwxrrRu3qGCR3bZW2MmztpPpcIFzsVKdbYdrArhie4wdsfunKVBJaHhzLeHs6DNRn
+mNJBtg9LFES2+VQ5K2+NFBxcgc4/RUYtxWPfT+mZdDNFSgv+GLkx/HQaeyWDaaAKMJ12X9Y9qrF
cijIYwJmgM4b67K7VvSr9Cdmp3vLDgCqzM6d0rpJiAIx4ryZgvyYuQLpnL9lX5ZBDZ4wt5ibs0kW
iYt5hHnTW/jz1yf/DK57aLx3Oq8XAiSALDMyD4GpHxWKp7EKFWdnbuOYcF3oYB11IKsLQMihT/+M
+WrxJVxOkZHsm9xHnmthNkb+WkAkJkAPKGnwOZmWk6h2cqmFRb1AfFOGpoIzT1lPSPhq4SuLWjKL
QdmimwC53/nrPypkMQq1DjcPmscPhpRiFvIdeqorwm8VuWiIRnCFHE6Ima/RQthxs4URn/VgCJBU
qXm3nt0b7xIN0mMKdsWcK4Z+8Jqbxcobj1mn1woM7Obe6pQGOKlBh93/nEkNtvQ5G1jY36MyQORB
cvSQ8YtOVfTZJWVXDA1X86gKnXsvkGicxglYBPBpxf3pq/bWdkyLMyYPHt1uCgj7wSyAAl5JR3J4
QGwGhPaDxGT4fA9mcQN6bbYwlHJuZs7VeGxGhGXwTvQdNZst3VmhQL4r+j91MS3ju7jV5JWe1vXt
+/cfpMiNTGWUDqIDAaZz9tRQpvsUzzxl2KL0dMbvrK/qlusqfAzcXSbOdyzEgJnKHSpuE2CYV7+P
ywNhs93kZh50qwLCUnI8Xcq4M1QeRBEND4tvg0ksEG847XkstFk+TkRMuObIBgZUcHsmBRBkTzPj
LDm3QZsLu/CLfDov6xd3KthTrCv+OT1La08//lykLWm+6UlN5hJIZOfWH+0ENaaCCqpTHCdE2+0p
bGbQyVXVfFBZ7xomUBm3FXX+WnKENU3Wc7X6oO5HtHEOhynGfNhRwdvlbJwfFPsbRrBuIQkv6ILp
0Z2zP/q/LHPRpPYKPbwiw1/Li6z4dA56jqta3J5hivMtPjAxknw6piqGb4mx5wrop/RSPMQnkDM+
Ao9jON9tOBMQZneGLVBWMy5JBLvQjQXECGLX+NRoAlzh0Ku5EINrs7Sq+Hsk+iy3IGZ0QS1T3E+k
0BeLKR7rcV4AXVceAMMhc8pO7JB5jOzDBwsZE75xMbhfdnaTdEPHeU8354K4myLx/Uon9UB5CeM8
O2p0Gf/fs0QJsWrFsbhxevh5kBkYQUOJTm1aTMMiIWosuraAXsj4cS9PZ/LLMY8d/AfozKlGLt/P
HH8H4ANSU/MmchZXjl2CTsK4u4Z5JeI95JS+9tFYy8F//QfeqiPJYAC/MIpZLV4dWfK5+sLbzQX8
4gmsmQqPIevvpfXrab41ENHiU75qlOVzpegmPHAbmrxwE5VTZ/HOTYHO2S2An9DPbVFp0tWtlEFa
dxQn5cxnIi47etJL/tJ5M0t1EvBsg4NKLBCFFtD3vdiwD6cz9AS8WzVtIGabvC1/JJH6vJha7Qmh
zvPjj5ZH9wB5JEh721yFrvr9NqKoy7FIvimLBMp7/RDVWjvb7Aw7X0WU9ICc9SpUrrVWCsJnj2ze
7mdsW17gBHKmdq5p6fN2cwRlCzRk20GqxxoSJ+DUBSJeud3FWysMIBrDt0TFtWAA1dlfb6UQkKnP
SiaYFHldg1qcxEAIrpDm9ZxeTOi5PANZTBMOPPt5idXRVoZTytkUFBNRRgf7Xz3MfHIeewJvUsfM
kQ975VcsEC9cNMKvlk6Vgsz+gbbjwSJGYICC0gRbGOlek7zB3bB6sVVYtgwJ2PCwjYevDL5blp2v
Q67mNT5BZ9X1wwXa2If+nL3kJrhuR320uNKZkCSi2LrgBRTQ4SnXhHalvuBq1L6xNmegL9CR0x5Q
07mIo4KA7UpVk3gzZrVTtb9wPN5Gs5jepjusGtrs/Ne4RI+unnMJm4+1p3lUkf1m7KJG+818C6/c
jKSSxQoK0eLOQ8MPZcxYS+bp0c0jWtiWd/ap+Rby1T+btgZVK7t2Ev/FdMRUKm2pg6NVZMn2ELVL
i28nA7MOazrla48LxrJf/6hBkx6m6ypnNhVW0TEWMaNOEzntxDm5LS+QlmU7he2+h1G9oJVXpklY
fSdos4i/P3WAe23rJ/jqTuHtVTlQlxnTvLpux0sRUh5kkPk4NwcQZVoPew2pFceKq7oMO8YKyTKU
6zJKJSiluMX4bT4zk39OvnTB14y0kBA5WADaJDddexhwOD8yiQ4FsCeGPYzX2w9GDPuCfPZ9EWCG
YVoXBa5dofhkEges5WAyXmXWjMi4ySxFRVinSWRuCp/jTmSYmKbyYG4N+rwYgfqAdUzdMLphgJ0y
l9mq4CVFBK/WvByncyxtPDAXIteZI9gf3Gbb70nK0Li29DCWwVOhfd65JR16kY1linEkpdpmxdcq
UzervHiGIcXoChLD/Bjl+ihypphhhVtyy4I1tXBUF0jdsH4XodB3P5USDiPBlbz5wXVvvfJ5+0cU
NqPpR5DFkUcqHqlelPYQRXuj2ipcCF7ZG0fFfKm6rT5bFt2qVfpENaspyFZEvyiqexVZSrmUtPbT
7e8X3R62jrMhpPiJFkOMx5a0qfYviy0ZHty1TYaq88IA7O9uZpGcheout66DKND1hHhQADUirGvI
KpNWc4WhfXbFjQNvp+0n/Nm7M1mowWMc9HCne5o2hIikLPXckysXMgmJkLoKHYaYVz4WCbF6zcu9
jgbr7q9YofhJU9/4/X8nUqiIUdi+QjkIP2Ean92Y42KyaSlAJWdGI5wkH6nrOeqC6ZAmDBUSpA6y
sACSNJ2Ws5fvjMUAxN5GiN4WpCI6KSV/40gUeiWmRZgz4vEX6MJ7YLmbFjKv1+LIgp6ICYImVDj2
kyh68PzsDUUGElcqub3he2LEspSDXz3zdLjyCgLaIi5KZu+gs2mEqnaBFBARaxPh0MOTjnzGVi9L
wjpoWY+Iv7iaWyg7+HyArPhl6Zyi6cmGIgbkpbkMuYY92UXo1lpDF31sLuEQVmZUzFq2oPISZftj
gmPyT6xqoe65m8QMmgotKkrbC5kTJS2yvi/cG5kysU7eprUm5qu7OU/Kv3Wwsz8CmuzVNfG5lBCG
o4krt4ekZi28ynu5MK+9oYBseLNEN1bXI0/ffaNccjkwgB34cHq2gbG3bXQLRu37rtT/jrj694hc
lSoluWqSRl+n+jkIznH0UmWFWr6f73C9FdDHxaRlezkToHqIQrI32xFzmteK5+Jzv1UeLrNF4zRi
BHsqIASTPAVa6t/wy9/mBKieQ4k2Y9UIa2PCnah0HSSFJlC9D0DY79D/YT6l20+voXqDxQTd0Xu9
CCB5zVCS9jx7886RREqE/e5hfl4R1jxLehSpn33E2l+Gd5QP52GUcafmqCefBCJNl9+etnzyoqB3
hmp3gjBwDu/XK3H+KD1aCjUgjI/Wf1crI7ZPNwzTpRlTGyTpmPUNXP5BSuZBZJrbkHpUJDzkYSIk
vvk49ThQ1hJDFVrnQGrzFuW1VA7cD/Fe2778U3LrsAmT1ngPV5WeUxnWiKhvYaVGtdAGO7O1Td58
upLr9OcN6WGrtRUawLbTbif4QfPkY8TXlD2/oorMykBBqr0iWhi5Q74pCCN23fvN+qwra/jT0oHI
Bo9uSuUwKMhwFRwuyUO7bJOH/ejMteLHG4wEO/NI+lV5rHv+xqa1XpWIhiRx6X1fcRciJZeWNtmB
5V9iDFFyqtEiVGdhywHmxFN2L1RW2LUXgswfwGoprt/tB+vbBHdk63Jn+3ln+yae9KJxmQzUBaFi
/uVZbZk2svk6z6CJS5xPsMv/GS4lJwMATbgUs9Mj9SFdg8bJZFHPNdBQeZc2sPPhsKyq3j6XCONX
8t7G9VDsUQOEAFHvlqw/nL9FPK0MULTRDO4hw+0qWF1RsVziLloW2OVzSe7hxV7BZjwQ6Jk0DV4f
HyZK840uU9oCRaznTvrBFfQSfYpl6psPI4ZZMPWgLH5iwVh5REzWoIV/Jk+9lwjhT68nd/1CEF6Q
arKntNbZtCNFPVjQPcVg2TPmI3WZyS3pVR04Elx5Eg1jkjQV6k+aiFvDNpnfeRfvm2K7hq1Lqjil
ebQKvYocAavo+GzDJuKP8QA8Ln3VV3xIAsIMn1ooutrAvwn9XRuYShC7BUH613fjG67jyFQ4VYla
a+PSQzZsbaC4o1gkyVXTW7UEixP7EdU3fdjgWJfRHs6qZgLlwo38w/4W/UUythSHhMThNcn4wxcr
jITB3XYnPrhXStABVuOH0IgYowx04ZJq45Aw2Zd4clNz49MFhNHvcLhkqo7iCK1x1xeu5IpB3i7J
CHCy63tKr3Wfea1IBb9chPSve8KhVkPelo034xjOGQ95uJ8789ons/Ew+1jQVn1hAOuEFEAYjzuF
QAazz1bkQKgTu1ByQQa7NpRCIqkuj2E6ULoX/V56Fq0HZbxpzMrnAkCDDLEIvYUyZh8vtF4LQMgv
M38ZSAWQSqgutI0qpF+6Nt7TBai5/+HLPphZaeI4Zr9aul7hn/FtEenfS9mxfmB2kmkS4GHwKODy
3w7Gt97RKIuGLE8Wb0VzuP4nQgI7c6VYYUnanBZ9v5hCsWh1pxa2iTSLaODNgS2vcPB0une/ic5v
E/pBhWX4cxri5Oueaou3CmB2PtdYwKOMwM6Wh5HjszT8SukgrZjHMF0Pq4pf3+IkU1ejRmATh8oY
ggpg3VmsNndzzVA/EVyZosop9Kd0Qf1ZT2+Ig1fxZ23NhF0BH4p+QzPt74BZU1BHYTfzpQdc4PnY
PNLT5wAoWZ7zfzLrT+7SYNwXnDRG1fj5BQYvdkcuwNxVW/peiJ/L+kFkXDHR8JH4Fa6z/Gz2Vi7W
R2eCUhAE597ObnYAz0kfvk+3NbQ/z88WHW+qe+/ZmjzC5LU0A8RlUkUzBbZQywhwCJg033q/u1X9
1N2B15Mbh9/lnIjDl3ZMqh3oJf3lEKquH5dmdFbbN0/nRGfyNxCkHWTI6tOJoHaVtIMLDnk3HFWo
eeGjJhKn/XitD37UKYmAmP/Dn0VteLd1SHh2tcTdM+LD8oUafFPY+XJU2zquUKcrcgpEs43ymbyE
68y9L3KXgo0zDbaaM5DYTv0El959onz4NOiHrR1KdWEuTgi4c9kn5xomsI0MAUhFxE/tJpXHAGnx
HLM+4OyXzBMcdPBfUFZiEotQ294anvfS+laggpiRDPwiX0J+uNRKY9iEmFVwI2B+MT4gvfQvIZeI
XF0KGjtNkCmJxClK7Lyhe7i+xiLXvIi9WqSSJAUBgzlUpuWeha/yNjIfPC/Ha44PjD/yTKWTX5Y1
+a2t7Xd8Xqs92crH941OAEUjkwzZC6TeyNpvNzscENwbejU2Nt47eLzcvrJoKV2IusdVtVdBZMIH
NhGO8hwNADha/YkyTh/eO2ThRUHQ/7uk5Ik1CeSbas68T6vADWvDBk6fSU+1edB7h1DBk8du7zvO
Nurb6qKO4r5I7ZM0lGRSb1EkZ1KXcVHgHnpsD+aGSLswGayFtOqhfY358dW7iaTzlDyST9aHYt6v
7geHR+E7rDtDQ2JrDkFFs76NeVmFr8ONObV47e23+gUy/+LmXdv+nExJZFM6R0izV2efUIAeKMHG
BrGEEfS4akqH9CgbVq6UfAw4I7h3fJPLhqMHUqYWO7eYbiR7PHT7/UlbZckdLWgYRof508O8Sb/K
oni+wCxnwoOR7kHZxwuOF33/6HvrjuxnGUU+KW6oMI7tPmQjMFObCv0+6EtUiihiy2nbvsrq0Mn5
g8y+VIyV35CCLUvolmDBnq1AkdiKQRcMju0LeaxUT8V3x0318vlso3Zrj8HhqnQU7kINrKD5lfeN
5ae0nAyx2NeKkOro4gNTRHIsRjUxFfH3jhnuNNjqNdSaM1GEQlOR9I6JNvXHl6Ii8ArJualrWzGU
ncot1yOsZwdHjc4ov5h/y0Ic0+pD95OqoNTdT554cYU8pPX53LkNxjab4QQGtApBeBT87TXxsHEw
h01nlOU5u4k5ESHIov3HtUbZZmr4Lo23/bffj0z1D0iaCGFuecjvrFxaKHtzZ0VDns+m2wvb99Ly
5m047Ol5Z2hycHQq6tv6Dd4SmaYy1ul1Om3+3I0P/IrZ/m9diKtyXe2NciGq4rUpPMhlVuciSPDl
iYGWQAJWkRL0Ujl9I0AyDe9J/hQauF41g9Ror8MrFADyROwFhihJkJTzfkELygQmsU76KJ8DzLiX
W+iDgtXhGpUGcgg5atvfhhkb8uARLv3klZK59dqo0lkZjIQQHZFs3cJexBwFoKZWFKjGwL3F7pxY
uBQUvP0s5SkNqzJZ62fq66ue/AgRTzdJUKCFKXsQJrdDYpz0i1YLZiW8e9/FYn0kkhFhZyp30pA3
B32avhkirufPCOK8f7zPlfdNwsamdQYXjkGkliLOtsLWEz3bh1rAYM6Yp4mSCq0YlJtabNJicL3e
uroGCfKIC+H46lswxvO5xmoVztAMWNQ/iunsmb8XK4bVDSOaxbDvtXuj2p2+gSzdMM9Ye8S23Wdu
R8qWkO8t8V8PiYP6dTJTLtmIDrGf+4oEZ/165OuyjH2tdT3XSkFEaeAmif6QUUs2OUwm3XAO5O1/
ZXbIHRNXHSEunfsjYwBpUoz9eTyGw+nrReF3Hf5Yw622MkV0/jYnNGud29Tmq26BX6fiNuJK4uAc
8W9EebX5x/gGgyMe++aTDmCKwo4Wr/s4fwlFkLsWRHXerKcM9wAR5QV6OwKz7lA9iTMcVsikVUlw
0hHnwj8DFtPqvNypcYFUCMoQaV9WsvZ42Iou+rf4C3KVzmav5Mc5WZKcvy8y+Z8y39zs0hPKh25P
gH0bB2ZvXciOkvwTiBmkWhey9MlbdmNw7QI5znDNuhwxA762tZQijmYS2oQdc6r8aYZsskidq+eM
4cTPEVyNSpqDP9hiTMKiX0xLEnXVsyeUOK84GBFhkESY7kKR+npfroBhpbtSgqks/6BXUIVlI+1J
PWrPZEGx9pPiYPGd35ibWxb0kY93cjdzkA3A9zp0Yyf/99r6SZP6eW9PRZaOgC6TDjkv+H0SsbE9
2vc8+nsUfhCtra72w8yPh1A/T7FxXnQ6ZOgnq7o8RX5s1tyV37CBbgSmJT1Ey0ce8w/964nbUj/T
pomPhax4rUDxaCf+5qxIVLkMhiA0vK1lYzdG17Cobpe2rdnssbFd4IarFjIZPgIFW5+skAje33gr
aQfg4nLkqbb4T1jcY63fyCyUMh+dbD26ANp5++Ri7jJF5KENJ9DQZNBrg962bMUmt56nLFiY0avv
BUIC4cI5mVG+kOxvo1gMpnAEwSBXl/fgf3CHZu/AhA/fa4Uov95N5t0JE23ZdZBDwjHJch/9ndnQ
kmLEj+vKKLKOS5KEuc4yUSqVQoUSWyhH4fMhD2YBWwwjM1IzdmierfWUjC69nnxgAusY73TdoNUy
bw2lXbCLe7uzm3sfF+4NqTeFt2hbKv/aZbyKxjLlRFqwqPlFzp+KEw2T3M3Z8pSA7Z5Ksc7QpFw4
xzRSSbprwiB3r1/ejzg8fhDlKV9MtcbicK8keQvMIsATcu2wtajNxHKA+GOc5G0uGvh0gQ0PQ9++
gHRleFWnjtBlc46ZzYG/CWv0NkF/x0DrHNz9JrI+oF16ppZqo1nX74eiyPDCGl3RD48wIKKP5kbw
VzyP1eEptBsmZXdrzS2hebHnaav5/NvQ/npcQrYWqStfC6H1eWVjJafdyCOfJ1yxE9hnrmJP2u1j
k2fTgvdqwrTTaJDftXw5kkSD3yIN6pmt1lQNmIEvFTrBui1iQfISTQ7lcMDMGody8MXgHVdO4LIL
GjeoZn/EDNCZ64Qew4yewuHX+hsr8z5jK565Oz8lahdO39wlwgGkhU3nUup9ydRBxstxQfl0lVe3
ViJOaaxD03Qc9vR+i0feCQxdR8w2uMhN6zJwInFDM9GDd2Dte0Tx5nzlz12cCGeGouFMYBf0lixn
pYaN5V+j/6xj1tMPBH2IIQeYdNiTMIrema9v5gL6X/6MmO5xM/L9GCau+Bbo3NRjF8lfq9QcO5rr
49Osh85O4ur8FCNPbBedyIdlwENY/cmHJc9ocnoB8eebzaaoNzaIMr2/eRrWsSgJBHEa87VUc52k
0+OEXB14IKlxs367FWYspBysKayrZG43QdjGtlYswFrG+E94RCnLZKw6heSPuDBRyTSXik6lq+Pb
h4W45oi/tsTtEH85+rEqe8Kx9NHjM35irUpojtrk/3QA//+KHH4MsHgTi/Gbz5fWwxsPSAgK/Wr1
mWCEOdyiU5AS5YGSzwD8zvM/zUQPzAj5+WsmCxr4FYu9PHK45ePY1b9ZojdPuAYPhhJeKaEJMLXi
n+2ZvJkwPFloy2pZy5rzVBzkIqv9wLp/PeyUa+k4pXQTkxwZirXy7oBo8dmR0OzuDacTKeZxNgFa
mJCVIn9xfhlgPGRf23Tpb5RqSkK1UBzSl6hHeE5ijlCLm67//kr+fAZSNwL6cjEQG+gU8ceFYfSU
SGwvnr0c5Cz5fUD2pL6cwaPoW0KVEc3z8p3xCajqyS5wtlv0lgcNz7EyTcXbg0Mx6U3vtqhblnen
br+VLgVWs+9wxoLbAth0Kx6fFhXjcwX6QxYwKHBovvfr0qvbQgLyhYcdF1WSTwKQ6G3GOb47tJAH
9Rv5bDxL9vJvagfw0tBRvnxgrS1HLRAAbybbO1735Lwq2Qnr6OdN6V6lsvrqUrFxsz97CcNxNE2/
V1CKbgw8fv2AGOwVpdUV9iInp79p1rPCEW9vm8KjZKl8nnaiPqUm7xBBieJ0SMCOJO0drHO8YWls
/UbM2ClbinJE1yXhTpMYMo7sgNdceOTNDGg8nwNV8Ybzu9/AsBhD98hTAasgloWYnvWPt3EGJ+Go
vRM9bpdVgL4mqcLWq47vI5EKr/jwV+ChWytlramiQ02V92yTIfj3i1W+s4P39t+UDEYlakXjVKsf
K5YjxUOIM/Ao6TaYGBoYtDqj1pZknNB4HaIYR5n1wLJvh6zksp4V5JMUcciCsRRa7AHRiR0IrOwN
odn6sdS+WvvXuMgJwfft/WLzGFjGWC3Re+lV9GPSGHwv25XOHGfaO4GxqdMxoi3lonUJmGWochb5
1Vyi5RR349z8jJoIt3D/fFuEpwpXR/cN83VlbRHs9CpVUjH0nerVS+gWO5WqspY0HV4wWfWlBkHP
3jZmmCc15cmsMB9jpb7CM98oc/HMV/bwSvXfQI7vYMn33EffroUWklp+dZ0jZGOXn6oQycv2vCnf
8BlHJPtdF9mUrbnBmoEuaekcVpeUvRKRTTBxfM2cOYunrB0ZHDdCILAQwHIQGCD+TJPQezkCw3EO
0QmTYzsEWcYs9tdBWd0GTQB2IHQdGWGmjQN5WLdwOzcP4JIZa31wrVQVAUKvY/ec+q+PuQ+SRG6t
CnF7jHwJhAESwHBrLeU5mctaXzSTSjP6SSat8MoY+OrEHhpDvz5AuIXCZHkZzY2guHm1osWJwRS1
Io0SKpCT9+GkoeIPaelPtESp18htYzG4GDwIvtmiKcMcwCnrPwRmp4qbLr9o4dmyjPP1FWXpmUKT
okTab8FWfOlI/YR7LiPwjgDH/hJc+OoX1vw4Yfm5DLlqac9LePRmoQQ8ZgddwPppa0zO9JduuPQ2
9U1ieoPkcgZBKRhKXGG05U3XfMh8VVMDo8cta3BjaE9A0fWecueKzQe+rjG3Yiy49iia2IePN7x0
bXFH3IEKc497Aq66LXu9WA0vLb/kUp070372nnU7Hf5J8WjN8kxioIiFFEKJPs5Myoej4XP0gnAB
IXp8dTUQ3WDVat72+NLhpJXGir98ErsxaCV1ktomY6hfBaszZ+RuDGlY5kahRe5zQ4nXw06KvtJp
bqJRn+litPWiM5oolWmVIeG5TxYFraBlGAJ5xoyUyAnfC7svRD+MdzS8+OLBcIQfvIw+TZYApieE
qToRzl8FbY36FY3Pplpg5IO/sy7/OxTkP1Vvh2nB/EL+cFHkPV4V2Y2yel1ZruQBzH12oHsvfO9k
whrwpjVNPtlzNNB5bbcnTE4RRwdMCW3+OA4Q6ec7MW3dLHD3l89tTDPDKcEjKOoWne1C7po8exR8
Ww8V0lMDkyqNGHlAPYAf5G2Dv6z7q550vEsRfJR/JBjWdfEEXnHTz0xm27cIpwEIaJuG/IZUZWs3
NJPD3Xf3XKHM7xVyhuX8BW6y/dX2Hz0ExUEl59hWimJZG7OfIA+WNu0LMesJl/ZX3k9/oMR6Q7mn
ZYOdtTEF08xJbBNyfTrtMEIKMUVZGl0wiG9SZKGbcczZVZKNtF+j7Z1SURR/A1H2SnQYxshSCthU
FZtxkTNI/tObRo0pOrpDAy4f6UQTa6cNejQsUUyjYfql8bMPKkEZrgWW0ecJsL0w4i12qwi8pLDB
h2CLkSPrn6j0+PqRrsBxJ1cbiWywhVK0KEmLBEPeMtda7im47mL2QFb2FFY/4lGwG0RRQcFsG9+f
sJIAm9/ITyMR+J2V3cuRpRBzu52AWV2DNaQdnMuYBsYUm7gTO0CxsuF8TwnY0TygDkQnegPURCz5
IvSKJuFVcJrEcfr/YQequANXkFE5uIpbszJgGFRRNrcR/6AHplC8hUJ//5qtXcyTx6YKORKbgSPM
QQbC23AjMOPlcqwznd+OQiDAQT4FmT0vBY7ch8vsAmkUc+2KV5uvmi9Avs+hp4VjaPjZpNFZCpwv
bG+es5eU6w4Dpy3b7khfsOJlv+thsAXPiZm1wkk1fxt/tiV+tRUin44IQh6yD3w/MkGebnDjlYk1
0clWM2PnwR4vf+A0JFRypqH/8+avpB956I3zEhdTDA10KHCi9X6D+VmO3JLeO9qJRJec+jupaGZX
B4l745PX2JPRW2Nfbtc9fQpQMcmlhkh2tMELVTlotU/0TG/SQ1KEXj/tmjC7SEU9IjahSLLbrsui
vhQVmbKBGL4ar9rGL9VqZ82ZshBWccmRg6HgBwlFajqz/HynmzphP0CTKheRTjNj4JJCaRP66mR4
NGYF2f14VDh4zMfaFIvcPZcMfFTT3jLrlnm00/n3YJnHAksRNzWBLanGKgb1JQp0TYuzuCpqwjjG
s/+/oYvKjxdB+AQeF0Nxtm0eJoo+tjWJ73bYBj22EbJqJwkeDrT72nlNMH+zoUavJgAwP8KnoXFN
H4hbPRs19tjSPON5VHQMg/6fHJsLC0j2OPLFLIrArNm+5F72r18h+uozA0AMiaYERC9xgdSyHxmc
JwlDs9NUVHiIWKipUNhLHkrBQ1sH8TYL9CZ+DQPTrCg/0oQppqQ4Lym03Yz9HOJrbHuMKJ6qpE2n
/KCk2GSudDc18kazZ+QfN2/+74QveFYKUKSesl9DTdQOEZOrUXnnkMffC7fjgJl2oF+TPesRQ/P1
NnPJR4vMDHRZX6n18aNpPgcywCwWKo7PsDlgR6QaPismpfRF1yhs8l4xhUl8644dd80/ArqyOPS8
lueutTTWwnWGvUCdUTgHrY/A8MCcyvHcj7HEtdzwH8puhml1fZyFX5jfYFZENKlYyWymWr07stt2
AtJ/0JMQM9Bw9ysT+Jyk7hknaS2hpg6SJty8oLPSOqJOgcpTgf99OEz7UnBBDcHAcdiy5I9uuAGN
aP+7Z3Z5KSEoTj9GpZ2ah0kv0YTabP2mnOtkghQkTg1j9F8wXELW/LyF5cMlaPHtlcj29/pp09hx
BPMR0LR10t1BJuU6jqZ/tUTN8MH2iCVWIQ/gAJMQxowO+qIdbwMdsh0W9tZSe+TgncjE0f7VUfJk
io63WM8ww0YBAqamFKHCCi6bsMa6z7b/DEvjNQLUX++Gppk7T1+FkzlPoEkIEckG5phBEibf5F3b
TupHNGRbZvrHAf2+bNFiHz5HQD6oQ3ABC1HY893Z+DVPv0EUAjk9jCoz1QFbDwqgFRAao90hqzJY
1jfy4JGIZuuhCIv5kN1CiKlw/UYD71O3TRNJ11Ti4A1RZEXohG9/1D0yvCVzvdje8yC+6NOlkJZ8
GtsLqzKJWH3Clqjg2f+fNHo2zx467kB4Ndmze+j38ceqOnselQXA3B/7gx4W5EO5nqp6Qbt+1uUR
NXfaCq/cjhkSuVsJhCyxPys54QnIHI/4nSa073M6NJMxOpwd2xQjEhWguxetPQ5szBJKegc3Gai6
kT1GevuyqL9RI0H4qM+qUDRokOnjxT4/wG2CmNuRoGP7mQTd/wfaeB7l7AnochPkhp9EdZr66VWC
H4ma2HSxirxZIUV4LhM6Rn/XI1EPruTBmpr35MnhKa2h6cFWVjSt7XyySjOtACGmcHSxlyIsvnwB
9r9YwO9fgD6W3uEI0NWOyI6XQv6H0GnKPiylTynd96ZcAl/Oumg48RcbRH1YCKCP5n8BUoVTD2J3
6Z3BqAQyOt3z+sm/3GcPtyZ9DrbLk2ylMMvf7IfAzGY9p23fHy3/WU6oX5r0Ne/jzeQMWdwSSUQI
ln+8F/VoJ6bG6e0EWoflcFGGpaLXSEjuxJcCiNSN9vyOx9wVkkidrySOgdnFL1El9SwMRFyB/bvP
VAsoLVjujXTdqIGfuhygpTUvFNNZJuEJ7IYv8gl0p8QhHJJ8GicV4MGWWsc2aFYxQ5Ot/wBuRHCF
av/lALECIjeicT/cNYC/iQ8rd3FXQbtqEIa22mbhm52oQFjOtaa3qTjB/t3nCiwDBklbVp+n78Ix
WaFUjSuC2QP/xgwS3TpFg4XvSIcAVJLp5Clra2vUFdM1CuwH4nwV8MbeEE6UpmlMzQemzmTU8h4C
i945p3k+Ag8HDWgtgDkrYV15ubMgYvuzE+jRkM0z31riNrWhKBFotiYNTvvAnIBY3lZm0rdn8MV9
Qc5YrMa77eGkss1J1TRmp/QurRNCCH/L4T9nXTdWXzRNSEps3QjgFDAE6o4LraZ7zsOhTlEtr6Yk
E7OQUdb1TkMmQaRCeuRzAkASDhe0Wyrc7+/t7h1UKBbmaxcZCXu2BruKvN43hL3XNrVzCGXzp0No
VaO52UQUykLGpeu8LoILLsd0LAfXv2FuzO3x9fvSq5XgdR3TJJfOe8sIkfV0pIuDo8Ql88EwyOYV
owCc4lBUDMXLtq6boRlcynhZI3v4tgwvY09jGYwRsoI3Y8ktNtpHRi2Z/iw3RxZty2rd7iN41G77
hpnqiU1kyToPEH9Cy0BC9Ip/8LKGcXQfqyb+46+8cmvaDRng7dae97WM58lTB+B2dt8Ei551E+OO
O+9Q3ciKV6ijPxbLg80uhOpQkJBE0jzOYNnuzjdtwDJ46JjZ3Qi5QWie5cyevjpEjpnNHUeViL0Q
Q5/QFWMawSjubXpoTEhl+BRNc2mp1fRLMX3fs9uT6gzT8PUb9WBMWZfsbJC1y65SWJlcmAqAx3JU
OZIDQ7uPaAZITUVfIGR7N2nzcSx1vz/RW+ZXObiixqgtpm5c4/DbpSWg1oRUSefWBbTkeLLGZNZe
qd2lZu764jtJzq9HcU2ooEsO4oE9uYzj1TBU4MYkj4QkPUUQgXZfdClrvZ5wZyaRlXM8jjFKfiCf
Sojp6zWbbtZTCmtB5cERwMMMY7SsZwApQsPaydr2AQPJ8ELZJkNN5aMRKk8dcDJt8xl4SHkTleug
sorL1S6PzEnamDqmJ/8m9zPUW0sPR7AHVtb+KdPJk9UbSw47XVCC03UNsdV6cbzRu8sgrty2Yo3P
MsvBM2exYPgg/NrNrVXXRM4zIVlfllt2ykMgeSnCaHT9mCOQ4FSB1ZCUZ+faEg7CdWMk0FrcWLMv
lED59vFTckLk3iFw1B4P2UKvPqEY5FyWZKVuj+AN1cEaH9skdt5/rK/8tUWRTif7YGB/4aGcV6mI
bLlzWWXFNUh1dlNwqRwVAcGNs/19OkTqRyhRkxhb5sgtP65VA6E8pIcXPguGn0CNUW1PY7Kvr6ub
V3ynG9MiSvtyJOqTsUQbZsGZ9UjucXsuAFQoXce/1pnvUvSbB1vB6Vo+tBVozX5c0xHreE5IWfvH
okrQ1NA7I2XZpEyFL5Df1pLC3KqOXDxMZk3gnGs5PYiA59DOlqNJkaKa8L2lDccRb7BBSK8lt1v1
leLGZ/up34Tg9wCA8rnuf43qcjjuSXR78/F9tX8zv/opHL/0ueJGZASpfBl54Gx+ySlCA4IgY1aK
pPDmhuW0WK5BtQ5cyLSH6Zkm9QsIpnd/S2BXzzyFpqAiX550JQt1+2DCyyXl1R2rJJ/Cvw5aosSQ
T1zWp93cc0lQUM4zrHcoQdWnhxnmqQ5lw1gH40MUwBfg2NnSxC0fyTlwqAFgzgBhRHS9aqjIyV9n
iMW3MMohiKZKpCK/hvd0iSQx8owsKbbfeF1egpzFtftQH1tMxlFVxvkLkq8hX8LQj3IfCWK6LGGp
LKlDcZhv8gSFVjFXGbzXNLOPNf6llqzdhqOLxz64PyskmLJrQz1QyFz9xXFN7csc+SaPkficE0wN
/PgQcdmSIjX/HuJXz1g4AnYZHz8poCYlUUd2mM9CrRQJ3av4D07ME4mWau0nzraAItKaXH4ca5PI
+kiuZ3t9tE/y7rJExkiGlhb8e0Olo4cyVzCUFnMv9ccq3oNYjfWc3naoCfZPL2rkVJ+epsTnLg8Q
0zUUd+wVnB5nLdeUYVo9mPgjeOq1heDPG6Tv6W+oB3BHfdkUOPwjEzQYR+OZ26ZR/Gi3WysQ8C1e
sRQya9qz9Rqr8OjqZf6fN8AcSDJAVKokZMlffVLsU3M7fVsQF5Y5kNTW9DiR1K1/dkq2etNajXbE
jW1CKe3BYQUwCjwBv+jaTBGoWG7UBFYuR+ovW4iQgJLTvadjyIRDtKuYnzdDRob1yQVcBLDTyIXo
WQ2lPatkOsQE3q0+KRHQFhavLpgJBS47lugS9wxwyYg/1xvBbkwGH1cY8rDvCMTG0EJrYZ0nW46y
fQVbactx1dzARcTTglJ0SW3E7DjnxFjk618fRFYPkbwYojmsz/Z5WfB0If3fqRexZ0tUKrhlLQZ6
MY+8XGwXVZi88xp3fe5ZAC5lROBnh5WAFA44gmN+kJFtMteEJym+htbJo2W8QWNmcefix+pIgiXB
+TBftKepTeilas1Nkmxy6KLmm6dONooqNYxlX5XJDd1aisBR+j1aFZRdMsgYxYA9K5TD7tWqw/De
x0I0iOxb2p/DewinnUqIXuT/YFOn8VtYaOR94TV8k8SS0wBFR315MW41T1ekCSSUccIiJYnvTwV5
ivqYFMJ8RwmErh2f6V+9x8ERwCgcIWYtzwNwGLluixJX+E/g5385T8eVptNlAWbtoL39ZWkmngSP
bF/6M68e0kY0VcEiSTCt2s/HSwOvOpTQl/ewd2ivsoXbTfBu0cg6DhibaHWbCXLr85osF+XvOLTe
rrkeu045xaBwocLKZZy5oq/uNo8lCnYDBf+Qnob2XmWPA+Qx3aNQGqAlAS0WSKkHI3kJEM08vNSC
QmL4Z/1dR9b9VD9Uw70p5suyGWzKbhRHLt2k1T7ErgEqZ+nmgAYgzYvxgD4ebMe14TPwncZwQpxT
o2wEX8MWNUQb/qnKxvOx/RjyZulWAzyj1nNUGXjlZHG/X+I34a34XJVSneS2X8cIK1KdMvW/j8bW
h1GVi85JYKHMEpB/rRTUg+1vF/7RBRzVfkyCpWiXI0WWjsW5aea2TpcJuvMkV4K3mS4cuJfImFsm
nIuxz5vbCQ2d08/Y3AcAaVur9DYcSOt0BxMe/hBYL9QgNUkYZvHkm96FoCNQu346uobV172RFFEB
yEfXqWh7D+TNYFl5qP8i5/CIjhy08SD++qqOFiRafLNGA5IzFiVp3O7JIcax0xzQZ6MTGMZa60Wj
BAZBhGxkPfms2/TE1eOFUDeShO/Fp8UiEU/g0i5wNFIeHHiDe0zdK19W/9XQBe8eaEq/iGC0Tkm2
EqYP16FjF+z4b/4io9r8Q/jXkO3v5wpApIHF1puANtrSD8Gf2pG66YLFKqYa/kxh+G0Ih83ZGzKa
nPqSWRpQeJ0achhu95S9WOY7j3fJeS43Cr4PZIKgw3y/exdj+afIsMSqx9+L92annIiuu/T6Jwwa
ticHyTE1HFgdCrIBRUlVtj6HHVKW43ol0fYPErBojiom7sE+CGyunj1gO0/dmbTibKHnuUuulFXg
GqAQ4MfYLO4681hNGMn3A3Pd+WKcHyJeJ2iSqHw8tr3m2MhPBqoGCs78gniwPtmf2TS9/qaeygCq
xO7xYl+IJRA869uNiY3CQTP72r5vWQEUJXLi3t1QCq3jLIGIfofAj2HYr4TlzQbrorSjwJeos0R8
nZgE4t0MPr5DR/WaFNYPdHR9m7dDNzlrSG/Mm+hcZ/KfiXuso89D5bumGlLo5MPL5EQxrg+kjYrA
vumH7tgtRmAA2da9gYFn4eLFk670Ny97RmRj3FDOpE3xXpr38/T2UGT/9FcoP5Ptk5nrUbmjFjIs
YDiU6Ex6BzVoLky3O1zVdqkYiBp9Tn3MJ34NluOc9znbMgyL5FQ4y8TbE3ApQW2rOfWBMNG5/YQV
ls71NoL6daFZ8oV+X1hY/6aMGtD+idajvHZQ7vduiaEHu65tyIU8IKsn3/ovkSNG6SaVkaN0PQB3
Yxn/2mAGPQrrREAMQplyyNWwAdViSzk/moGFYlagQdcK53ZBWcxTDiejPVb2WH9OItnew3tMiP8z
K9vtGFJo1/MCdBCU7Hjy1vEQ/b1BPfIhUEv/dr+UnPyUbWXQGSvOCBdq8zLeZ9+dIzPZ0r0dqxgY
Bs8jvC2pUESyiQ6hCWvaMHz+fll4UQFN4IiC/EX0mCUSgCFPus7r66VQcNykLmwrijuZNNJX8z3G
KWsTPvNOBQCLTPqMV/73MQ3xPQ+vwIzcahi5eUOy3W5EWCLmycDlOpRKmvZBBLLBg7XaQDaKX1wc
bnbg4jcwUgibqaqzI82YInXKhoECLmduuWFq1Dh08wDprf8Ps+7hvkd7mebJEOO3CIo3DAEz2AMe
8To8b+hvHg/qe+eKbr4KKyuoHXbEEvftuXSyfPYUlgPzuby+l4T1ZluXVCNq17tITNBdTaDZYbCJ
TOUZOUuWjfdoQptenFbpPDrsgBuTpmMD7czUyqD9PtzWXILNEvk2fh8qUkb7y5/Ps3EaEMz9P94Y
1wS3S/i4u6hgAarvLEU855hBUxxf75yyNbwlQ/b4mXvF2xnzvEzh1N8HhnkAMcPWCAGZV0y6/2+v
2XfHAeljRiskBH/rexhmetFzOL51hnrcyOnfqjlJoRPPuslvgr/0H7b/On4yA3Q2D+Y4JRXJKDUn
4FAd4kW0p4wrXLf1GQUz24jcJRzZSft/UGFwLBC41KVX07SdVV+8GIMJYLzLQevGXY54KFTU/CSQ
PxJfsc4MvjfXClOUKvkplfB5hXSzrw2oL7UnIlwMe6GaxYl6OoPo+e+bqzpusveOGx4qo+pNAYWg
GPd4ScbHARlQo67LRn4aI6tbQgz9w5T6i0P6Nfq0IjTd4b3ufRI2eZr0IaUtULrU3zID/OXxavxg
mNsTPphvDgMyiNm9DwlTZ2CZ7VH0DgIW7Szcnc7KXnudhSdNudEO8X6sgMEhU7YueaK9Bp0GgFJY
curwMLwH1r5hvDjyOIZ9V1R7dUEQ+0E5D02g6NSE+wmPK1wdy08QTIK7vC+h3PJlGYJCoPHByHbp
DX3sY6I/aPUPP2MLMJH3LMAe14huOln3exxevzwCgecFnsn7zPiXiRINMwuqHwlDRg1h9k8aiWvh
vmMTjwewuAPWEjd0VBkAcNLdOw6sn5jothkVXIKfWBpoQ4IcYsqB/RGHCwCdhLF9KD1B4zM5e85s
W7TVWQsLG5F9TPjemWFweGe3rtnJYkZSHg4F2xRBSMkB5RGyAYxoKyodt0vVdPmz6IddG5u4DoYs
s4iNSAAf+fdNzJLgwVVlXrPL7PsidTvUU6N6DgYmOqbyIGzHvG5ff+4HaNLWntz6NITYLkfolrzU
WbHCuEM+na93D5Sw7ljlQwidwBK9esNyyJbPSMlYOm4kKUaelSpRnPmueHr4a6qIV1ElPj/8b7ZA
EMWaVgBRXPbwayXIgf9E61HfdE62iVvAKrjyJjTOa277Y5FvFmDE2lIht5lHg4v3rsZj+OfEGhro
W5fklxAOcwO3dcG5r0inyyknoJBphSB0LBF+q5JShF6x5BhrSksYorfJPha5YARt3JY+kguTr3mg
CaI0qWLSbvWQSGExfrdTNqtXEkcoh2LMQH82DmpzCncdZhuDZp0uZYfHIQzsolr5pEMTu6TIlGQ+
DiMjgalsOkTDv/+XLVB4JBeO6+epCKrIE41tpdyBq0FYnlYRUUmWspNIw0LG40BlBzO9fa1onFI/
IGiiHVvnr50RcT/fVEeyZvrN0/V9rlR3V04cud0sT0GOkmVkWdTXax4ohJxGzU8QrydSorccM58o
VvcbJ5T5Arf2F4Lu2R8TUERNhRqyYhvE6Szv4OjUkOqWs3a/4+07d3GO6Q493uzT8cDnDnO/l3/c
buQwUHrMPyQO764IQ799CIZWw+JFdzZEIdH2IyhdJqyCXA9GuurGcSoUdDUjLrbxZDm1rzxMVCSO
fqHdPrnBthx5Q56Iy2DmS1fQ6o2bvzZYthKspCjRKa0Iv0X1gfY5BYIPihS4tl21qCjt3CJGaU3z
OYdSEk28DP09ozdwgqo/0MF5mWaAHjaqpQpmbQAxnf2A5W6PH4/Iu9EosOZRGU2IwVCQ9rkTAfUG
3He5llrCAytZqe9mMNvBednqdbnghID9HBMMTbKj2DgpQibx7+n21pmakHMVe17Z8Eoc0Z2PGjl2
94cxdbF/WFbHrFVgGxoNq4AmcN6+olEvi4Kawh8f9mlKJS4ecITGLkMCSMaUdVVYz8hLHi9f3PBK
w8VK4cq6ZVdoGKWbH5S9c6lfQrYHf3Pb1pa4PrfSzPnLVsgzBkTnzsnSVfHgqvh8+N6gI4OiEuwl
gIMgppsTcyKdfNMTIEIIfJw6HusttNmWc3fMN54r2a1UpG45NAivmY1fQtKDIe5ccZcVXX1BbWyW
FvFOnoOpPxypTHwnOtmltyuYQNwr9vN8BtInplDAQL4uv04yJ1fbWzC2Wlk0njg6TuVCV4qd/VdY
TYLEy7vec7BFXYm1985YpXVEdlPGHeVxIVa1iDhbltDGeX95nkEbR3Gkmu8rbs07eVrAF6Dmem9V
jovp/iFiTxbdbeZAjWO8Q3q/xHIhF3BkjOPKqduSmfpSUPz1bkaKD59gppIfo1jQoWRm4NAY2WRX
6MmkOipqp3mYoRjYZ2dWaKTMb5IeR43ahriwpa1lR1eqGQ1VSVtZKOJZPzXD8uTEguFnKlNLzjfr
Cy1TzetxXX/rPSLyXU9OZGDXZ171H+wTdaREYnNAtEPTykU7XQQBuQyVELqTsiAF4rSFthMoadZO
X50a7QVxoaG+MphE6HuV6E1S5ZtpfwS+Fe2f1rIioXxwBQelwz2iaGZnhpb3ocWhoEuhk4LG1jhb
kXt9P0g36lYUcVzaN+X/ayVhFpZt3AkKrYUd488Ko2kgVrbg/dVZwRPR+Qmrd0xjozRLqSKeCHsG
5KmJcRT8G4fPLZRhigaURF5gHd9LMieR0f8tPxUK9bnN7p6oBM5HBcRRifSMnMPjF+mgpiYbfd7D
qTEJIzAPsVwjs9aELRVnXA8B346zxhvR/GXUnD2ob4MTIthfVvhz9SguBGmTkjFBzerIAe6ENP0R
hIRWR1kYckCfAj+2z+Rhn+faNEOjq4wzndZv5b/QOJ+JAHcphS6V0IT/pUw4LfXAghyMGWyqhBdh
qATwBZq+R6NbbG90cs8hI3IMrMg1H9El69+HDRABnkEZn5/Ld5+CyhNJEGgkoffAXrsA9kS0YaTa
NYCt4wEjPyDcazool+eKc53yhPL+h9pJxr/+iCBCVhg8YWf5KKX8uUkzcsqdslzhV6BeevNfgNJZ
PYiarV1WS1WOA98/G0OMmjYZvoIAkjU8tAFr0vARuzGFNvFy3ckozEVw1x1kxKlp/gETInDfLyEg
uzqqG6uD2Bev/UrLRwGsOwSOxapfzfsFf/riI3NgKFJeo7QhzEQBd86ZvEfXB7+Ctu9UjFVB+X5T
b3HcCaCPonVgFTkPXP45y1O66w4Xl3Eq9EFUHfLRdsdjvx4CK3YEWa59aM7xajap1rynOzFtZHgC
4JYeFvM6Rr/SxjgA1OF6a7NgeLtRMy2R41im5GiRljrAYUN9D3FkYlfenEeIxi+CnH0RRjVJRA9z
fklEGmr4IzUAPNGsLHTyNbK5sYt+85UHxLo7wlvgzwXC9slWaGBV3Vhtl7htg0CpY/kQGxlESTSw
Xre0Txa5ZMN8wJLmE7rA5UfQrlryDABbKk0eKzmBy0SrUFKQSPb4yr4XiKdFMqzdTgIyCLErcrlY
g9CZjfOnPKULKgGs4ubg59pbfsLTC69Mnk2dInfLCpHhXaEreekxbggH79GRXNR3WOpjBzFM1BC/
J5Lahi0FKPVPSWyp0UmR1NXAch4pXh0uB4gVUOll8rjRMzZvNBQtM0OyDQd0FHFxE6zLaJ3AxIpC
ZRuPQgd2jm7jS/BaHIUJrvbtXCou5Wb8b4pSt6/xfGM87rtr3W8yMxC8z6fxaJx4cXuv3QrcKgh0
fHt8xVt3xrbL2ix1+x384uRYtTGlCiFXzCFTxEElDyHwe1zVSLrtv70+Y1YZW0xDGzFYDfdMEKIn
vmsJF1X/CDpIzEQ11oSFUEhAlS9tJ+4NefAVE1DHbu+Hmbjz6e+fCElOxMuB/+QdQWmZVLkWuy/X
Yx2w57aFjxy3OtSG2fkdNrVvpt9Ir7JSJCqbmfz0V1kbo14nP9Pgwbpp4/v9ugGppe8hMUf3qKwF
9SfNP4Bn1kt+hqv97NDZ5iEgGcLrbv6CNzbp/WvL5CKJ9pqV9ANKqpfYqPMOmQH00KF8kdtbl/EJ
OjZH+IQXSt3k3CkNx9saBOizNxX0B13eituGAVC9KM/FsCPoPdRn1ekxoa34+hu6XAAIWjEztiHg
swpDT823dQ8qaryo2t/3me21akiCUKl2dnJDLAegyvijMsbJY12pqy7tZ8HhusHfehDS3GtZUh6j
4UBiyEdVOT+B+Zm5eM1Hib8mhfvwvoCClDC3+avxAYMqRxH8ouAgh8uEeqHeODFueD8WG5/JF4Os
NleMZtPwRsCtpieDZzmOxDmxVBADrX31JcEJqQ996jqY3cEjmsAoOFofIrloTjyJJrzHXwhTUJ+S
nYpAZqprZ6fXRTiaRSbe4zcXZFyIbMIx7j30TjJyyNfhoRiagRE+QZQtnV6PKtG+5rzQuMS0GWKg
wTEiGcp0BBGKVQmcQPS37UVKf5KTQe6OAfjGLJWSeVisO9bU73D9f2iQwnWf9fhB/ogL0UfV8ATt
g3ETjenpIIAi+S0UokYH/AoOtyCXsVVCts9T6j20C9+IWP5IjZgz1Qjq6BybOWWJl1ed7uh+5Npc
PYq15SxhBP7aCaiEw1bxSlowEeq7b1dEPDtjCbiW7gfAOD8M++8Xh22Y0+TH4peOxaWj9ZNwXqKQ
a4KqQ8qDhYJitgQsKzSU+1imttsag69AzRVeUcyYuzzBQGqGoMvYx23MkOdyNmt+KUFKt0zowyxG
WhF4GF36X6KqyI+ARJUHKxS/kQtz+WAK7WF6asjFe86YyeeICYQnKhnklceWtPpCI7gIs0hVCBN6
nnQcKF8X//mnU2GUDuZyI6d2EscBPCWojsotYjbGGKOqqBvq5xAgroa4oVy/7n0UwJLHRkulDktx
0rIc0hLVEmPyUZmCVLqkhWfcEXZ+MGZK4n97TRdSx5hu4Mv20YhZE6iKMjbDsZmzYZKoFadDO2Ch
cmIs6O/NL9byo5cm8ecdvi4rah4DjoY7f2buZXCT8pOacX1ybHXTlZZ4hoD3t9S6W3pEtrTgibD0
5Oi31IzJfnQ6AMpKFsxhXuXFFbRagVPwO2Of10GQMrGs0ZIpZqkgebe/PATOas3tU71MUkVAIOSI
Xn9wMhcKWZBNf8gJReyFgW2J0UWf9igPJlrQVpzZdDn2BSsgotp4jkZupVNFpKIJPJlaaa3F0N8D
pWj6sDpj0ymxPF2qnPQoqx3ULvgawER+PG9s307ugQDmwBiZVSHd/a2OEDpPjDbBnwBjCuBqwCfT
8uei/GaMZGct75Re9IAsY3Nq8YYvCq7r0jQtXT4PhDt31jcLD5/L/ESFiHYGFwvEN3D8EpW4kUsT
g81B5VZesGK1RvjYHs0oYvcaM2/nBqClzOLiXS2K80HLLetJPsS9Vpzj5T8Zf/vSO8PsOy97mipL
MderBRq4P81VUrv3OQsG0l2kQzgXQf6q5dqiHZUqNm4uI70hPMCLDqGO4+750iBQ1QzeHyB9GMkd
7GqgVTFUcZSP9eLz8JhPzgfR5xjXkmPloRIuA6TpP5HgmXRit48rnbb8y4/TIUH0n0b/WSKxWOSU
nsJtYijXeY8T3Ty3Uv55nw9o5vjepWN/RxIu4TYpe/diEXmC/Rl6B38PYdg0iRoLEmW7blDPE94n
XcUFsbZLl6IsXbt+qmhYoEpovtVDfCKVlgjZpJge6bqDhWSE6ZGu3zs9c6XiHt+CvJjXylQ7uMYs
q5zjgSq+icFnq+oHA/qj5IixUcPgu1gsQz5t4DbkwEU2b35zDehlErqYxLSeLurkUp5ksLdK67Lv
Edi4zq464uSa5gVHetkW+jLnKAX9UIyYTOXgD/uOHxv+KTcMsQDALywfcEpEnbH7+8PIIx5kXIaD
WVgtiOjDhw1AY/i7+hr8bU1XiQjbzuNiudAiByPY9948P2bic9DDNN6jqNnbkKt3ukMjefCohhOf
jvjZCmEHBkUPQxR9SULRbOPVAgjHOYLxRZ/wm6OsLBc63jzp6r79jfhqYyp9aB0FgaQEBNe4xflc
4CI4VQ7dcuiQVMpVB0IBnSILgMIeGwq8iBuodxuOQFAvoUAtN8cqMKFDTi9YE4h68Y6/tRNDYHDO
Sp/Vv4zaDEB/Yr4d+mEWUG2gQutc2XvkDyr9wHm9P5g/LY0D3v+Tpni5Ah5hPT8+57AhVAzFscbg
pGJykv+cuvNN4gEucQP+CbocPY0h5hRzyw3wVG9BYqngIY9jYEOfDy6s01dlrwaDD5rtU52brjxX
EDbLMMBQMFMeP/LqZcQJiig7XyPdl8wi4SaHUCMC3iUslQSxuWAwJCqkUq2bzvTcVZfx1f5aBjis
k4j9fPyNCsOgmY0h+YMtL7kfH9wRF3N06+0RpjJFRdEXQL4LVa/5tnd4h6cFXUH+BYr2vDCZ73qC
DmznAJNtIzoCb3DDDFBikjQg4wEH4HRnJtr9EzylGfqaPkgXpIdJ6Cd/hMF0PxPruiGwp8Vft8C1
y95RFTlUj2jtK6tJBEyo+iEcne5Q3K0wELAD+RnqthBT3cv0BTw13Y6ZaD9QwXYuWBIkYbz0WDC+
p75f2jlnm9erSc/XuV6u27Di7xjG
`protect end_protected
