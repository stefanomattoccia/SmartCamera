`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fbDaBFHIKh52nacy9jMzYCMG1Qperci1BNhS3a905yYf8AeecKbmEQtlgupMzzq2Jx4PoYceu5dv
l8wFyM1beA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Utdt03S3Lz7i7p6dw60Xpdtn/qfD30vK9yxGkNw8JA+BhbYYcx2eoy6xX3s4i04F8mu4ZXW2yaRZ
QiRt02sJxlPynHgxFzZFQmLJ7VAzJcFAktOKXhWNwj9wLoAbrMTsjoWkKcK0jFv8BD3HlVd+njar
EYmkdb69Iz7LBFGQbpM=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4PT6F7RUlC6ulkKy8EHrmmm//6hC9n04KErb4TQM3+Jh/QcJmRo2+sfuzcdUkdDM5tVLyoL1zas1
82QYOJGjRNqJG3/ONBtWFb1AfoD+7KRaeqKM0ekCCP8CRxqTvi4BLAj7qKoZYocNy+9GHsu6grZb
IcibNZIQIW4p5GlkwaM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oXpOej2si6vfmCwhxT9L2hA9y+uHvnEYR0CqR0g9lpI35C5OC1domnau9GAI8KKsKod2cMYkrO7N
p7BfJt68O4gx3HP2fnTtvSGQPi4hCU4JENf3ea0gZptV6Uug73DvcxlphHzEsfQvNDytZPzCDl9i
TYJRC3+nNJ17CrUuAjQw5TNZ5CEr0ab9sR5vNiV83iixbHVzhRlMWTba+N49pyQq7xLXTuw7KA6M
WgaNEcIO3uhOCpLBhnmF51V4crqXW3jbuHGHRN41+3s4eLXkbwxVGgIXBKdxNE2911IrZwlBIEVI
fGVkj/T3llHvdFKE2enmfnBtG67VsqyqSxxLDg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p20y5FqSsxVqxQaw6mFQUmXW0btKlvrXp4sdgMO5NU7I0yS2G7wUu4HdQz9aEDl9Vee8yKfezePv
lKk2Xic9pdtgGsPnB+DEqIub2ViadwY4ObLTLleVBZgq2zcbDjSiOGkRKMcizquTL5/BcxMdOLUu
02Bsp3MFcDoxOYy8ciUkJiA5G1i57Yyiw9rCwr2Ta5+Yyi6RtbWM3lm8yQGLM4PubCTG8tkHfClF
WpFYFE54lHbdMNH+GNHfUIWynJ4avx4pyymRgZ/1Csh+uO1sG+rm9LtQ+fJIOKsR4UqptvUtNx5+
dQXdpnubb2XNE13HIgKarr4vtrXwnd05n+buJQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lqz0XM1L5SrgMWZTZt3KjAQO8hxce+rwEG22w1QNMgpWvLZsg6hKjbPLKUTF5//u48F5En6+esxI
KuJ8xEbRiHqjxj2/3FhHbQyfyNDY71VV8lk2FNFJtZH2lFJGOj9F80zlm3kmvhwdLSnrMDCci0t+
sOA1BiYTZJvdy5WvwhrJhOJ8uGLujb5oc2C8InL0jxeZPku4c4GpPs4ClG4Vaqujl1YuTHw9nwgT
2VoUpAezNIeVLFOBUSIkShA4NcbLqfGZPQcX1fNAoKz/yN4NE9vB82uLm5W3b2B2JjJoX2c1QSoK
msqvphRnK2MpZEXP0f4zktg/gfscI47gPQFk4w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4624)
`protect data_block
nyGWB5qqpYafdnMqNNuNaX38zRIJB7dihSsoEz6FlQ18U1vgYbX9ZBqf5y2oU4YJnnNki2fw5Jbt
qg3zKrwToUNVCCZwjtd1i8ucG7ljvES5I1GQbcostnOVXPMFuwaX6ksVCbKLEYdR+EFfkw/e9wIQ
3pFVJdn3x4yfPMknRlm8Nbhz/7d271mwaQgKpHXWH6uKy6tPwbg3+zMNyv9bF2kMm8ygicjmWBk5
p5Lc5PKj1by6/W0ZDw4YTVRyHfIfxeeiHkcgmgzs0j92a2y9qKgfjN1qJ8nmndwB9cKsOdCqCTSF
SuMaWBSvJQ9aM84wnXu19KJC3E3o0HlHFI1fZWuqzx9JtPFprzGc8yiXkjz5Bxp6zGN6LwHgAHQ8
JHAKH+vqv8FcijzV/qbC4qjVz3RHsbth++bDO992wATnN747lqfoqV0kXDB6PxaqGuv7X/PRLpMJ
FgTmqLKv0OATxyKSBlqRBFlLh3szr2MWR0YVrKfeQspz7AUdxKceqmwEyBlUsLxOLvbz9JzYx57R
NW7em1/+ECNFVeNVut7AXMNipfbwcuDBc2xzs01bmrp87/1Ut2mC4JPehPxmh9e3mYpSQI5+I7W0
XSH3DTXBtAgL8Dxvp3oCVKmRoj8JsE1BuZu9AmdSYhbdhwOwU21y6SRVFqQ5jemfHsR2s/MGrLvV
2PGNf/WCJOgyZv0GMhZ9Uc5dHZBGEsPKLAQ7GJylVyjB3xscDeZ2JZIq77plauXHnZNMkOiV3irt
biO34d/yn/bVJoKJ8iJcAESxThzGnL+LnbkQiPzV2LkSayVemfvYoN4spsrYL00ph9pWGmh3R+g3
+fjzGKO3AsaXVD95rDg/DFuCg0f9WsD/wjgNK1h1UrA8zpXHn0EKbT9KChUXL/uhwAMAG1AXyIJs
vuU6kQQazz2QNbf3W1d1l3xEQ9f+s3oi5khDdunvUBcm0sLzmXxUU80SwEq+9ZHvxE+qYqvi+w2a
QEqZB1ntkkHePBjwBJ+5Q6MZZXWIjyODSvEo9A1pp0zlnQBNpS5d/FUsQaCmWSzCxocI9D/VSP+N
TIMLhciPoGyA6h7Jj4bW50JXGo/J/9ofsvEXJ9jJuemi2wpONja+FeoYZA5PrE31BPDv4L19XniP
TrbB7OtdmNPOTz5ywGRO0srW+MRVnE4heZ2qNb/j38hZpbdpPZqS4UMNr9LrANL3CnmjsTLVx4nN
v09q8gbMwT6nHCQu8pRBA7/QGa4h/3EO1NtYRMlchopJt1/HJLvO3JOIRjXWtu0Qc6kQRzzbRv4l
Kp0/FbkiU4kuCdpw1w8EUsrgezDjUEg81m1/lm+BXnqoGiVrOVlySsnW4wiwjsFoJDgljDCgdHVj
U8pvD25ScLXckw4ZD+coZka5Rn4IiZCi6D4At1k6g0O7/Fk1LvDdKdR0mKY+njAXgoK3iccKjbYd
XWF079JCFZHXCAh68qJ0oab1uXimJO805taSeNYlXki5sgNCL2CXWqCCT7K39PePP7QVe4Nzoaac
3hpi/uZ4z1iNT8RXa4Ovv0uCTjSZlqAlAIHnICgBNaInqTTJ1dBWOLIZaR+ObrvVUSZTHiPDcAAG
g/SEkXtUCL9ixBup8SKY2pRnzinnXXuZIRueaskQ/lR57VSYYZ2j1oN9tXEyGRQq0lNAWjGTdQSV
JWrZtqdOCSO9cYQGOWCWbVvZSV2BhBtf8T0gi7osNrLSjvuakSNuaUUvbfrdkodpwiZyv2haeMSQ
UHn34S9OL8VBQFjJlANBWq5pDMf2MrEi0/k8cnqGU6o0CLtA3RCWNesBXc2RLucX6tkWxJNqzZ7c
s1iwgiywcEEM4oUeFuCt6iXAXohl1xIiq/jMbiXyFD6iiJrovqxVSTOkDdr+xcRu2Feu5py4UQh1
pvwtaA3b9gW7VX3cti2fc//nyVr1sbf4EpDrBrE1mXHOJbX0O9gNhhQsuFzH7UOPHqsVNm+r05xU
yBsfsVTIIYStRDpsFpuoW2PpZMqMVvo7WfKhh0lBVziIWdOPajMSutUpbqTCl6ptpgKbl4Z2FjUU
72A5HqyEHv0sDJGJT6oF6GlS2ffbDjM8aE+aHebY2HLoMDuevXcjx5/0TXsVcs8qSJzDkqWyrLDd
76Qdn+2o0tp3Xw42n03WB+wdX+vuVHf6SVK9acRLMKO/uX8i+EtL2xwdYVmF92cyCeyUEa799e80
PFP64/ttbMQrLtZss9WVm1rCi/+n4TrhGd07dAI8WUJekBcOsgorpheGPrTfPgtXBsGbW9Un92kB
NymfB8G5ECY8H+N0wWM8WVh0Y77PQvrWTTiMYMiNhenYeNuGRN+NrgABSSqRpOTUZFyHXhzFYgD0
wF5aSaLuwlksfmlExRWmkD5u8W8MbxLOWW1TCZWaAtjBh8if3kxCBFAM2CU3NRe7AoThfZPbuUmo
hKxb0OruvVJFfoevufvPZ6HC4bwTfozb6hSMoa81jqMmFPirYqLN3CqF7g1ZYANclWfzeu0+5U12
xepl1TlamMzMKQlkYdyHX4bbogjxtt1rJHA2zzbn2/WmPCvv+kZ4cVICcMcqtf691q1fiyjJtTnl
QaXsL0DQEZLK4UOiTH5rDw+YVRR8eLpEtj+pv6GRxvFFI3sonpiDqYUO+Pjdq8ja3LWbv0kuVETT
TSux3eE3agnKnEj0bRzuYhhc5/abP0IrfAv7vr+h0pC8J3XwZVOL0orNrJk/SQUhBHPZiGd0rrjH
BqsF10QAsCzEzorDRTtJhEQUKh5rKnnbQ21+XEWWPVZNGYZOWFLiTb7DgEKeshbnFdpUSqtVKCl3
dMOnDrYt62jNT/swyltmEILOpQRWiCa/3eVGzOpQ3vC5aGzX1XJfi8JcG6ARhy7CfXnSP2I1DDwV
COLScXZzNw61v0Vbj/n0lPlHif5JXrewfvz9oqDOnbmnZp6InAAWUAk+soi52vIg5qkOc/KHzu/o
x+QCYuNFWgiMjKN/biH7in1toKfftDmB2c6oYqkD8fGEHUewIzwa21xO456yWlMPONZSwQj5Bd3O
mOouHBPo6owsG3A4yWmANYR+KSYGLK8nRxO5DheDURnaT7xb4tiA71lcLYC+/T8Cjv6yHNbroii0
2M+3pOKZfTnRIgfHeCE/QckKrrgepJPrjmyf7DawphnZR2w34V6nrlbFpXw4NF+2gC0CvBR8sqDc
CPLSBeukEmiHXABE9T4m4f16dGvWoAb+w0+rnQ7J6xcxHSZxMqED3j/fLB2LkcnT0bqVX1vmcdLu
w/v1xEFJBu/iXlQqejqFEG4e48qKnNm2m8gb6/YUwXncdo9fflQmyW7ZYZb7wpyvwa3LIBNqEXZq
RNWqXYI6M5mgzX0f5WwiWZBiY1NScGTNC4hn36skVw0ohIu6OnY20hFm9ImLmB7KYnikrTsX945a
0hMFjysIXoIZIIlw6YvFKKspcOuebNSpKv7lPYBkfU13QkqZ93mj9QrRNYn2pGMBjmzkNB5ihs71
+hwwculU8Dp23DRQXjBsa4+oAKMDOeQSN5Fks+4uIHsVAGg+w7s/Lu3ipD5EE5mET1GDkN/Bsc4T
qrs0pke+Ih7o3LVOWsuuiX8F6hFzPYSiIq/I5Ei8yvERLwSre4gEazhXMW1iXAgt3uX1x6cExQFD
GM1E0OHISlxYyMQpQ2y8KtAqSnTHLGizwjkO8dC5YOxtexkbNUPlEU01CXjCm3eNAn5Cvt6AXxpv
7kqdrrvYtNUFBCcobRLJNoWg2RYXNIDVaXtYkJ8yrc8Rl+2YiaObZIR8fvfPehx9BhyM6WMvvL8Y
R8+UFhiWAuSlMnjeVbzZo4JXE9g7spaXy6ypohf+u4HZKwR4bYXRd7/c1eP0RrMuEI056Sq8gJ3x
wqf04VHZJXdP4n/EsqmY8yD4Dtu/88nQTh+AFgFElq6mHcV+BOPHppTkR6/8qlFuVrSw+cdV8WEA
WsV+3/F9Foce6lYf3wAHHJjU7IOb8sVY5Ef+M6ZzX3mLXXzlowUkHct+e6zVTus7JN26vl97T+xl
pesK9wgRQliJR0x1x9OPBcYKDaFOLLbzdIXCfi9QjI14rAjSA3aVzf+JzDP0Y22aJX0izfxr6Rax
zyU7eeXr+XWZj3uosd74aHg4AmgSCqpLi3tmAA2DiSjOnOnpqlyKjfqi3RFbHLQVW8cZaVeY8q+x
4T6t34JqIbcz9OghgW2ninEg52UCUvFYInooCy2oTUnFP0fJ9LxyhYXkbpe212IBfCagyXTP5Rup
H1d5Ses4T1TcGpB6Df0dguzP9Y8Zug4MqH9csEp1rl7P8vzcMWC+vkHx3CUPX2Lox0yZWaLb/12N
M/Uba0xc2QuaRTdjP3QZTa/nz/4KTtAc4KTlAio+KNPjtiPnuO6Ylk2BiHaP14L+VT/MW8g7O4iX
IRJCkjJSv9dlEG0yvLXWsgkfTr2Ka5a1FReZiILFNTLaokZdr1TtDtIADh/cfSx11b4s/m7m/J8Q
vQmxXB+k8OgvZ6Nxzi4J4CEpwLEN/UmkdNeRxAK6s+m+QLu5LUnFC74GEx1rQNoOG8EE4tWxuvS3
LHHODSgYVNfJqnrtstyIFtEKynGixYAX8qG0QQ3tJvOR4ya7wEdvxnHLcK01/AFaJDmNvPiuN4fO
Q+tALpRIdSeldDEt41NI+smi136XHSuumaLeQAlvnrOnjkh6jDfJxFOZuRUWQGQOGE1CzM0RyvMP
ZUQidGUv3kdos+uEa3ahhRC2wBK5WL0sIYLjPEtAmRj9q10UIME/H7LvC1PO4vkdsenmi4b3Cg5C
Cvk2o3vfUYGOF6tSHuDkMMmjtXLociT4cvIDOtn3neVAghOj0uNt0WtUckyrISK2pdfAjzq3bfrs
0Xzc1vTuz1mIUz5m2+uIqaCX3gQzPb0xeRzXbYAWgLqEbCks0Lh6kUqzcCR6+pdRJG2VP0gWRgyR
dacNXeDZcRNd+GC1SQh4UH3uUzhgZAY0TdMkCCcn3RTRI8UVEEvgSRi2p/CxiCI7uG6BPPizIfY5
iNpixeuXn79SwW8POR08/3NHoRUlH8+q6UErACotQ2EMw7CRGE1X6VksUemxCSBKXvvMKkWBuJxo
fGweuLJMs/OZNtCVD3XsJ6LWlx+8/PeFPbe5a3tn943vbJrUCIm67YL/GIbrelQ3HHOhQzf+XWS0
iYz3Z+5Q+g5pB4HN9DClQFcBtwXIXNgmt2EPSFSrR2ZUCzm6XccpFUC10T7Z9n7UycXjS6XoHY9+
OeyyxjRyrgGhX+bfieEPmuEX/dTl6CSW4Sn4VNWMeVu/qbmpkpQaWmOBRy7zOLEAzMswdHlqGG0U
KaEH2zypBw4kkzCb757BNOoqpk1hEq+ROAIfc+4ukTnWrEMOG1iSAtH0IJQTlabGJTO8XawKZ7K1
Cp7BSKZRLQtYSmgEcfXcIFcXxjSh709A35vfjBbwArw+LlZwOdgA3vIAt7AHtTa2MsevuGO951SF
2OSNsatOcJJuaHOBQONx9vyrVtRfWNwSrnTZbYMFERiPQ6XrxOLJ9uGUWuYOM2J91A2j43ylAqBG
r4aUVDb24JymDKkvWyRaeTExpbmm85NhdiEzNxuac4dB2M91o/VMmlBtJ2Hu5BX3Ycwrye+nJxre
yzmxURECUQ+t+XgvEVxQ2ZJXp6u3eoh9FrSWHXONuzjhHOFw9KOgWBhip7i+CMdlhGHUgBtDtDb1
BvDV5bb6K/Y9cNqlFqDpg0e7ZE+bPPQS9cYwbY5SHkadVRQp4EkvdV87Ixk1PMKzDNJOUrrp5ZHB
z5bM+td3xv/ZShnJGsuciMCHx7L/oExu67Njqr0pd9wgJZrbS/vszabaRDFqxmpAJguWM+GOPkrc
4IpMy+q6NvImww5CyU6Rr2w0NP/AycI09UfbXXAxmQdZ0XK6CfN+G7ZhiKtjNBD24KdKFb16tVBv
rh5neRGc12FRik1cdWE3+KCpC2xjTGPkH2AYW6ZFxBCosIRlNPzyMumGmSrdIumjxap+Q/wdJfhp
v/TGXxJlw0vzViyVsyzoTWTUN5WDfZn6QPoa1fWCI9H2ngrhJIB61ZxuTPy0r5WoEM/HXRbhbpWQ
+Q7HK8fkZFE6XKwzE0qPmjubnIye1tno3fNpHQ+lBhoKtP/kmGZeVbn8l5Hq9U2K1X8b5QU0m0SU
dY6RM0kigA==
`protect end_protected
