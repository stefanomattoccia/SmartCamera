`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
A13f8tlz6UJG9JfCNcYl8NLUw8Tlctm35dCRvt/KCTpBFIuXlOawHL7sTHowWNnYPdFQNufThU2P
nq6r7CYRfg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oJAsCu5zl/OMFEQsA8TK81YQdELnJEDcFa6KQ0EHWxmJrxei82pUrFKy5/0YZah/J8433WTkuMYX
n4DxKRAShIrdY1X7G4VuvTy06p94vL5LjcHyEy4fxae5eyT8gPJ2ix4XQa8NTiv0ndfGQZyw3Nh2
G2fKlAI5x3f8zwZZQY8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wvBGFVtHjRF0sOMF1pCWFAGskoPwO7T2ijyj/eL3cj3Mn4RaSun2E2ii2aHguV5ZVFP65oRsiH5d
RuZPDUKAsxBDhHSsGkFSPIwX9KivlJTo2FZHlBDTlkfDQbn+a3fWxc1HcR9KUBo8QndFpzMmqgOV
oDGrjFRMryCx3hlDJdU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UMkVtIsRH0SCXq8LQlXc2SFapNVFtJ6lm3Wp55oPh2JHEa2eDcLuSNAMzka2zwzCEXltR/XJthW1
e74yTmf22SChtep5vBZ+ajUd7h2t8MuWnhQAMciHkyF4IkU7ju3JOoQFlih3FqDO3aUJPcamhd7Q
ccMUMAhIvZFp44NdLzl8HbXnE1qh9bi1m8qU8jMCKESUZ7pg4lNlsQjd+Goa1H9iXaLEv3OfHZuq
AS/RQip05I1DUFL5hACAmmneYHUVM5S4EEaO3aHf1jZ3r/piru3ZRDHXxDir2Y9zXiL2oDUfsV5l
w+Pp691O/rBEAjBLQdevDcp/mZn7axrfo7gedQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BizuB2M20zTA5t6lHKGfnJrucOUdZ0HEVkxiYzkxLH0WP9VZIREBo09OejVavblw0lBdoToGD/Dx
ZN2JWgxB3v9b0Oe7EvwN3oB8w0TKm0RoqDmuPV8JuY7RwxtxkHcrVvcjXuOt8j2BPe5Ix86NYRxZ
8RqRFVGNyOVCKZuaFMVHI+ktnNU/xi6ZGsd+L0PEmNWeJ+y+7ubRYuJBTcZK6n0e0Rv144/nsqdy
X+40+rhcynqZUh14Jaqxwmyc8eu2wmo21it2TUiXXzLiWf9C/rPTasxTNu6GgF2yKIv/qtG5zsH5
iEI5vhFnzG+RShh+IHFb+FdSgnifLxcvxMZyfQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WBEZpdyDr9NfPjFUCp37UUdIujNIa897wZZ58/x9eMPhksqlKdy3SYhoDdl4U5n1JXPWIonhbpyY
qfWTq0gV9NaH1PiTuV9w+nrQziNvPhnHnWOzNrltlMQ+uTbMRquXZffmAQGphp7ekw56wGNMIqvn
BRmPzqHv8wZfX/RCaFbjfXAJEmAF89kl5TL3IWnE72Kb9o1cSvFtKTxyRoh9m9E0ghJdkhnRh4Pm
wU/+pIGwon3nUS1E00edVC7apMYbKm+8akp/2UT8ovmuCYJtcE90yRZZaeiFNpLq2UTmaGHp3XHC
2ziTOAA9fjUjv2jhCi5RMA2D0eDmOlHleltm9Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7184)
`protect data_block
MlecvaOA8qYc6lt+j4Aa8epjicu27derY/ZWtIeq3FG5nRmO1LEw2yUXUZM729wjD+vJmZz4cXgQ
xw2X/yxstlNr2Shc9XpeWHw4o6ekomB1yHnpbBC4a6CJSCMYF2g+4S65F5QP8bQonaszAeUUlDGl
c7GHRNrKDDaxgrNowbi9qb+xuqrejZdTjbXN/U8IGSSlAApJWP1Z7q1e7+qK+UjiDIr34IT3uTPY
26ueLJKDcnoCgpHkHJpcac8yrwi+GwdJuoIFSPfC0MM2M37dZln8RZ33wR2AjXcHx7vHjQkjmrBE
7NZyvS+dzC4SxG6SxhLwOBn77L6Es1MuaVhR9wZDu68gfWLog08W/izRiF0vDwQK7GBo2W4bXiii
ncxFbJLFtIPj4VjLyM5EIHMuKTeMh+7SBKqZOh7s8SKmTnwhrpJtRF+lTolcgEo5Wv5AsLOfsAYB
s/LHUnGZa5ysEFLLlnUhNrK5ChzeoRjTrH9mSFnmPsApMrboDztrk5XVl+TPBINBnmjEDcP/hVvJ
OytFbuAQHhXrCPsAIdQigk+t1qBGzj0jZN6oKJzOI9yxlKT0r2UNXQN4Jz2mHIgSQtZjhd8B9r1x
jBU7ljwYts8yhGRRiyIG+PtzKQeeLw2m03nRID0xk/MMZTI1EHVDyqVRGZMDnLYHoCmIke0+LvQv
ntVwkgY4L3NVFv8BgRl1gZoYg8wm2xm7n+iacrxqAoO4BrKqC46SPTIgACERTeAoVgjOrP/8QpYg
2lNXAv+cq9TQmFbhfPfgvxXGLirrjxaC6sWD/cxDkpnYJ5aAtNST4sXBF2ew1oRCM8DDINzORLd8
rSVcYyTQCodL2Mz/cf8OS44KMtcmvg3qlogpxCar9KwLi5hwezEYw8pPxVAU0L+BJ8OIUmVsbw+S
rDeEZQbVBfcMIdLYQgsgia8wLVgXnCntijSTychLbBTR0FboLpyOo6nzJ1HwS1HARl7ydElrTpbo
g8qslk2DUN0EB2fdeWsORrpEkhxEpe2Hrn1Rqx5NrdjR7MQYqWRfLjpH41zkM8sry3nWArcMT2Xl
2MFIaL91I2nVCrU5WRJjvpRkKUvRqFeJxmLtsgb7tbKuRxXx8YBhjXsJpBgVPbogW2/sK9v0GD60
0JREDaxU2EunzCT/j7j+Iku9WkmKzg+N5U4LhuZp3TDUKh2rarf0DsdZAjDFefdz5BhX1j0igh75
cmsecukUh7+tSGXIhkiGFqPSHIJd+LzyKVj+4kEdMqf7usi4RrCxI+ApMKtiFJADLLylZxVbrGXU
7KbIA25vMe/X0TX3HfqA/z7CYf8IMUmBvydiknMG6qOLbvg6M0/iaTwbAf0iQFMbeRnF9wM7cGXq
SOvZxb7HE4yhBJk1BwtkqHhKPqiIOFFF/ap96XTjUmtLnElsmKM7PHIn6BovGa20QCLWoKdhUmr1
YY54VElWI30OWlTl09TKmd36qDO6h24IqZM6S/NNDF0RPhQioosKqm9DpFKpAAknZ+Imkf8E1h3g
NWGqy4+Lf9CMun841LNPNYKQfEE1hh+Qpm0ebbzA2nTEHqAXDM0+QKRQohLEaRwCGPbAKzPw3dUF
IEH0363cZ+/SQF33ksa5LC0hO9WxZ0aa/J4PufJsAvn0JVUMJ2saAMM7YrccdvzaRAekQ6syr4TB
bLaHUcf0/5gsRERc66UCzIJOcSprX1MrtF/QS8E3QT7GbDit7ndjETA5hRsJwcytJRp/FMVmxTmN
wnT4wFsqpzBo4nhdTWIDSdxc5BjFm3zYVT1+gCDIE2MvKE2MY0IJZYzRFuz4xS8ao25NSyyVO5YN
TUjJR81el6MhNsyVE68CfHAlAgC139uGvOk059FdPMFTNA95VBm+Dl/IudEpwMHyzEUyMTreURvs
dNvknYCS167GHKPiK+XE3OHlvNs9v8S4ZYJ4yCEta5rln5Q9R++k2YN78ScqgwCoOLV9vBqt488j
M42yCIAkBBOdxHzt+iQCoWhmbbWhb5tF/PboVdXTeSuYeNeJ/P1bKRsLOUn4Ou7JFFJKIEWcU4cw
gow6eD4C5R86OVeInVE5l2ypPgOJgIrem0Ne3XrwkXK89T3OzuQW5olMwFAPbW5kanUhNgifR7q9
H1zy4K/97C6uCLzva2IXi1DxmOVY6YUe2kyykoREtr+EGnS5F3AZUcKa/3e6UAELaZNqrwGBY305
n7dD4XJjB898sd8VZuDKLwKDn0I7n6gDilIAPKIO2fCPQto3TWfek77oP8LJ3+nPvp/U+xJndrGf
mtfKxhxA+MLRbbVgqlxPfrrFU25gqpRP7CNZGzEF911QBvetYOzG6KmdGsW33b8lgeEriABBFiDe
JtdmmIzxTOgXTgHMi+77QGthHp6cIp+TBJG+SE3Bd/HCBLHuJQTFs191jod2066tsu40TPPf+zHb
rgVgRPKhPSIxZnxlcmIksunqU72zsQtW9EGZbL5z065Jb7rKYd7UGTBrAHTCGstGyCAIHIPhpYQf
4alHA4cTUumwC7metD2o8o9xjZJ0YmrIvtpjhpa+Fx4zvZ7jgYJjHsRhQ2fbGzEaSz0Lkxq1KK6s
IUJoCMAr2vbpo+m75pAoFcZ13UTP2XCXbCvPuUYCWI8myvhLA3RTP9SNnr0JSvYuSD/4/2QY4fzl
uZpqYxm56Q04C4LdF1YuGfMJ0ZbZlGSvAlcMqalO9fIxR98jrtX1E/HFofxC9mWKVn6PpKXz9l+S
WD/wkz9Q9SZsIjQc9BLXXfEwsxhlR/8liU9Z6+2TvZKTzAA0kLYVXNqiDBg094uYwFoYFwZ0Tj0q
oEjh5oX07dz/6f4vnk0DgLwfEKgknrx7uaEUGeXr1bz2yuZb+IA5QY9ZDSI3gf4eE2cNbSXHUXJZ
z5CTrlB6wiwDvKL7fDWLJDF3y1iiEiZP0yGD9PN/H+m8aSACq1NVa3EFuoLI9s9LG7XRAzrI0HBb
a3mG1I7JUxWiwcFuAOPmP7EffAvebBazIk0ODQxaQdoNYxuTkNhzLD6Ti1iBKehe04LIB59MUDbB
fwwa/I+ooUKDPb/cXSCXOE1FYND1dGwNNQ5wQlyefk7Yg6epCiubd1m46Xxg3jHlNZ/R2LsijLnh
YHZbkjUHHKm0Tv8KWBdEBka9cdprK6k9meQ5LKtGeQi1n5toY0hs80niv79X13wG6HvFYsKoBxnx
poGUrWIM1mcv73WsjF7RU7Wc9LpYT777a3EsYZOPumpyWXTk5atQBXkth/2UFFOuG2GN2lneLdEs
bO2Xzj1NehriPN4nXiRHvuPtu/Z9gpX4XS0eFeBb8InTuJfHJfj4mQ8oQ59NOaxUfjYZPvw84o1e
dOgthDoxrfqzDinxDySmjCIUqGF/F+RoPahs8zmgFacH81sIYEdVBo7h61AtlT0oBzV5iXz74JkN
8KKXoGhP9nnOcoF8kQzKBMklKUCyqMBIEAJ2cGc3KgG6LXFeXGt/V1ENEQQMBULJD6Ec+KxIEFQA
09ChbRIaJjLwI58ld3wugjMXhh3MPxeAkcpS7zEnUUVah3gKtKb4qAuE7upIrdj2f2J/Z5jx3R/K
Orp9tphQiS8UfxOdnTEENsqK3LqCn31h3wqyq3aUpX0Msrocp0Di17wd9mUD61nzAgXw9/txkJrV
chNSM2k3DkQZmOAVfEAoHCRml7Ju5er3snmm09rswml2zHNiYJyTsr8PuMCTOCYK+dlTghDDj6/g
4e/WSomumlo63OWWFaf0QAy0G1OCu2wW27wMFp/ewo1SgIWTx9cDm+3kluysnWVxUXC6LvGfccm9
yajvkhpiTehJ8FhXZ/M4zVVvN3de3qi999VAQYo3y/LEE9yT9JkMZ1Ff6JKCINa0qCh3H0wSmRXD
h/ZBcF3T0Ma3nVT9cKStN7/GO3LSTHLWJf4T5u6DbjGC3lnTWSyO/bOS1N6Xw1of6JslsPLd0YE5
t2/Pxsstiil658W0V9b/XttgVY+1giNjVd1WkBbFPZ87RYQ/ZJNT46scZEJB7lysp2CfDkPcjiO8
qDCFVGBOvVQW5YC5h0bW5s+qPeJO+FyvxULPnL8zA+r8S1X3CG3LcNnbS+ykehiRe7onN3NIt/zr
wgkwZ+trQL/5s/dNs7ZZXwJ2nYjKuxCHZE9t4+PlHg0r/tulMDLA0o7Gbqp0lLdE0pZpr9daGva5
8LRthWGPKal/PYewmKtTaxUEwTS8GfetqtzU0hWf2+KjWgo/ALaXQ42W15QcgVkoxtUU+eiazCx+
w5yj0OcBYGonTj1B9ZSDgRxhqq08eILj60k/iZaQt7ZIDYEdsHK1/BFOGu9aMWSnh8wnUTCerqCp
WnibBv+DLJc4S1764puVpJQiPNMclYEkz5Ka+IchFUjynPVknTxB5KBQwLh0QXZVqZM6m3JKSRH6
mKmZQzvRHal86YR87TECyeITI34IlKOzS3CN3YmYOz5Izz1uRLg4gCvP+ewHDdQiPoIV/rSAdVRQ
tPetivjuqC/V+c4kx5XWHOTxbpOChLvfO/o3bjf5q8pbT2UNq7DzCEkcUnd/UGqM+uYZ8qcrjF7K
C7JzxuOA0Gd0cTdruA4PoKRXkSkA6GKe+q82lllzYoDc4Ry6V46yTQHZd+/EXqze/8ysSz31cYqv
IAp95V4Q8AgNWRFZf/RlLub5+uQm8Dz6KD5e1mvcXZZrt8uEyTPoPCjjdmZTNayg6SWeR15buLnt
l0CEDBYqJvgzsTHHZVTnIrnNkfpb1r6vtIJXHMXYWpsxvAxU7Tm15+glIhxerzCCw8Xvad+RKhJt
7XL8qivi93TG0kvZp44/XtsOWbOpfaIKipg3QyNjNvlWT+dJJGyCZKjXBlGRfQ9p+KRLHySms1od
SvrZbRvoOvVe8DKtd8xjoI1nZjyJ083cWIDKxutcrLa/uoaLiyTMZOddZOXMxtiohSpF0IqF7Dcg
hB5IJfVqaHMdhDDPpOVceJQYDCxAmr1YvXzeuGyAJhhnYJhpnPno+l3DKo32ZqvOs48rnQBQqCxl
e8l7QUOpr83Y7HqjSzhQdQY/h8Fh6zm6hHNc1CT0+ag/lPxoy6OR9oJRRArRNNjcdAIf+vfjwZbV
2fQK4iOhumqUTfE/TxWoAngBtntLsdxDJTmcx6yiGCCsEC9xY+YlWMHOiAAwofsv2eHAolFTpAOQ
s0YuarIeGkhack2MEkPr4ir8O9urdtTEU6qxqLr7hWT9at25gRxgICB4aMpiwoJJk9vWjeBdmhrw
llq7i6FyExP55gcJWP4g2nz7jjBHIPYpo6EPpJ42Odpf/t8GWJhIqCzs9p2b11hW16T9cewhzx1K
nU9A+qeS9fCS27I0YSJpPPD1EXXuBV57suAkJvKmFO/lwSyIZsuXBPSyptVtHap/NlJ9jsW1qsDA
bgwHIXokDVOK+NXBoeVFm4fPUuBvImBo2l+i03o6FMES97skJ9zV5n+sBsOLZj2xP5MLkkaEWgQi
BgO3V4dhKDnFQw5ZUvotvVO4dEVkHUbc6mMwvwQJJLV/LKKVb0/QBaTre1nY0j4gMemx8pGxHmJ0
P5hQMOi+KLa5bM9H8BusP/iZMaWYR/+szxsWrAfYBkkn1V66Vf8DXSx5ssAxeWmvB6ekhmmbF2Iw
Jk6UEpx6e7lyY7649HS6VNlcnmjZY4BRKdfpGx5Zc+6Ez5QdydJIZp5apTIoaH1/d/T++71MwN4f
tus6KLw8a+PUobQzcGC49jZKgdEe8lfDRVRZKJ/5u08K6O7AHkpjDVh2k1dgMJ0wTBalUoMFB8vq
haN5u9/AlOz2CGaNy1Ri0t2m4woeyd8nzoB2K4MXwDaq3aTmKmcKXNvBdA5tavw4S06vzvFZymJD
KSS8Tp2/hSJNyFJlWnxFO3hrbc8U0GjGemnwbCpn9dL5wEa23y1fF2fviSbXOkQ4+vWh4rsbRX7P
FGynTrYfb2i7cU8KtLLHuJIhvceg1d/pQfnjZz8IZrhM9MBDQfRnuuKokfvI6l1EJaelQSnFCXmW
UmijAvH1c3XIfWVa4J3mFdTerdzsh1JYFyVyoKhYzIe2+KjglvoYCA5ZEG0M59ezByISVklAO81a
DhKVMEhIvwwHth69oXR7r9V268GNTIwVXl0t+pLRGgKVmj/vDP+uPlwMKdfhA8JRYmXDuoRd/PNt
yeWSvZi3p0GRKcXa3EQFANSKQ4+HkCsDKJqvGyRedUeHEj/9O10QvLvwpT/OBNULD4N6pAK3dx7w
R88PsWcxaDEfFzOey4LAoRulT2cYT+ELBcD7dGM5Aas2F+Tn45JodZ3iAxtWSrlCZJTNh+WVtHWP
+J97oth753VFrnVoYaLs6wHqag2bK6ZTVoAVzWVXBdADv8ysIE7nUcJ1AeHYCiL2l/U8J+uapwFJ
N9V9HA9XYH4PHYRRfK3v/mvoXlQpNaGyBHXgcWzbKLTmoORE5qdrRDVUI+5fFWbng8EFrYANMBz1
LXxHWkIyYbb2h3qoFWetsShKTZ8eluI1imRgTVOCURQaVulhsEOhYKOUySVIMs0PDd/ttgzMUZrl
0NgUrPl7axPKLDDQtf9LMh5nbeKw06/R2ymZg5FkWoj2FSXkjCobY6rEnkS2cbhwz6+2D40B0MEH
hOuqaDALxo76WlBKBQ5M4gKCUh2WD7Rqqd2OdW9M0h2hfWihm5A8enBVmo0a0OMTz5IIK/ZV6Py4
1eRFtT/3Z2L7q9U7VYEkdtPC6tKNQvB9JpkjHgD2IJN3dLU0ImQqzxlxTR9YMLLgkREIuTIGly1I
wIgXXqEaTLBNqX2nN1ENl3DFMv8amE8JTnnmtTr4X2D+QacodpbIfPM12MoTsCv/cSAqczrQ4QYT
FD55KaUKS30KDpIeClJ7tm9U+y0q1Ow0LBUBddPan2O79i5LWfn622Mth7KrkJJyWeJKoRtn5ADF
EaScBqx/+wf29olLMpozm1CUIAPia1XhO3R+hsDADF04C2D+3TH6zV9KR+x0YoG10iAmP6JvJnkr
I/IFyLaqwQUu+rsi1HGfZrQ2Wb5duwwnX5mQvFwCt2t4lp3vT2HdOkjtnf8O1xXGG11FqxAKk4iD
R7P4vFC3eohs9l4gVqjNAbAXX2eqRtsKh1sb6LQA7qmbnBKHbx0kYC8tJlrYHScf+oNHAtMaMW7W
rT2Ug/nPts50fN8XSUEBm4SbYcANiWVlFpzddTbrH32cMVmflYSXPaonCEjY/PSwa/QQgyXEsw7/
hm0xe05ABNyQ6lXX3mVBiKiEaDKSA4JS3IuQGTvjxBWS5RaM813Ld9yFQP+2j3EMoT05GSgVElv2
aQuPEpVECPtkJdsx46GrVbgHuJqD+YTeAX/Std6Zw98RK+9ICbycE8KGKBzXvFb3X31zfcfRbzDh
I0+nXnP8l7r6NVV5UIvOJEB7n5B/sQmz30ZdpthCfRfI7Wh2CGeu1nURs7kAAR11npc5mzL99l4q
inEPhhbvzrGUjzMO+C2jw6zzIvsfm1v1Q6BabmEliVLraj0DAYYMgCIhDbx7AxwqhT1iBJbC7S8g
whltkNPfuTqXz/+RSqcEVg/vPllEIwqSriJz+8H3RmKLKVBMl2hCMzTikSzkRHewXB/IYk71dEhq
Qrx1MTelhHNltXbugjlErFUPIsSP84jpYF2BTHMxz8LG96mzG9Ae2vSAYYMjS0bLwtUB55brI3HP
nN2+0kzdPZzlfR8P2WFnraymWdi/ywHOnLS4JgLLZ+XGZUj27mp0qfBGff6GDWHjdvsIlqi6eLQe
jUllOYdud1s/UuJjrkcsF3UWnEaZ13209FAt6v+3Au0lJGAQkeHl1a/YIEgNoGkV66mWX0CrFZaJ
obb4kmTo6KXjGeAt/XAtKMMbhZ1e5Hn+2ST4kJIKXyCwboAGfTUcVUrrD7Xm1rp+pPNI9p3lmcjK
UJ28MN+LcdJK+rzKm3h07J6CKBB9j7vdxYuXapv3rHoSHmg27qW8GNipSe7cs/1URMGEVW/WZ9Ap
Z303enLfVFs4L17BWuwXOjhB0V8CfOdxhYntPEVbvq38adlc1dsy+NvpvH7JR51v5PvGZVuMSYWR
AExjcLBENw+3P1YGCoBvIzhMWIWOmk3ufoqync5/qnZarjXIaB6oeRWG5BcW7AvcJ+9tG2X0qlWk
xp28S8x7aQ0IBbMxuszfNTYsOpm49QUlWQMDueTlOSrMjQvuo37VHUgI4USweH8QKblzUnMpFrnj
ZMtqYwS68TAF/pooPsZ5snk07tazIZjpFRJxHadPab4ehXPBGOfXSGyiAj6bDx3em9+K+C23skST
xl+t+VsO+SytkBmML8TiYoDz+BldjHj5666C4q9CKQrwx4//Btkni/JwhwpEOKqkXfXtyCT7CzvI
dTeHGkTmq+80Yn9+NgQJvXO0gK6nRqsMWHliNexRY9o82eQHeeuJTb8fXw3XAFxuOd1v7Gs9pFJ4
m9KWBIXmAcWN2ZOyxRXma87HkgNF3K0ZUETfaLnqZoYzsswTMD1S+DdKV+MFY1mbmbcK6vVZxMnj
kuQP3yZFkYkoopUOpE4uPrfQbSjAgiXq7/8TSuEFiaJ/gPPy+TBpa8nO9814OTJnxk3ugjes3Jtr
p0r6yul1K5DyGHUSDTN39lLmPrFDXgug1LW3OOIYxd3wyhvnc5npri/k7ZMMySd3QG3loujnAoR5
L6yWJxiKGguFqR/vEAwfll/ApFaRrAFc6gV43ezJjfz5ba1dtCh94XN4pZJep3seruC29NHPhZgA
cNN7f7KA+0UxwXBg/TWYgEqjnYBQAdoLFt9n0ZyeN2PKqm689QznOeVRAQzvgnvCSHbKbni+jxyM
4kPwHAvn9XlnF0Xh7SeKgIA9qeUAq9w02HiOFqNPCXkaQvBHAJMBuVKNKjam5PFEjs7h1Un0vaVQ
JUXgkWgtLPV9XUvsTzyA00DrSZMO2aOTeqyiUtxEuRq0jYt+KzS8l8HjOibUjpPohjOARluTGpMA
uqUtWHD3ETqXDCSlrddYsB2/ynGwahTkPTgz61DsXrfV3eXPkmiMuXfMSKaQl1Wa7Kd9SUWC5H9h
6EKTqwzcPlAuZO4XNT9AXREN6wN/FtAGcfhcH9y5/0QEBAL65Y2b08yjF7kEkSCyl/zYKJRelfjN
QRf/YcICjlx83vVYtJpHz1o17bOlYprINZ6B/p8g5t3vPi4GUPmAtS+fMEQVcACKaZqMgUSLZu7l
joFBN4Fvn/LpxHR4/wfFSu2hni1ogCV9L2SoLOKXiNf2r1Zj12grWaKeOq1RUWlyT/s0Wp4ccmjp
yKvTCIAegtq9k9s1C+xjOGEWT+RGHO84alZ7a+O1zQXmx+OcgyMc32owiALsVSqfi+YcVV/fwipL
gYbLslxcqHw94GW7OliwtMlRyERM87/iwFclWKfLn502Bx9ahOPOnQd9rp94TMn1GT6EkMVqOmob
3t5OMnCgpMu9UWVS198X3/QnfmmqUFTXtgIfe7ceQc5PVivBWCBQoZQBZHimJfJNFNKE8AndpNpm
5WXkI5C0vwwhDmqelM2NwSXcQM6UFPwxzJNFeoM5/C4XTci1Ir34T5wEa7MTD4Km7pRxoTnzxnaI
KPY=
`protect end_protected
