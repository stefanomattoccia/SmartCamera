`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
P/t52Rab0MsHpvowZWB7JWID0gGmModaN/9c2I+JzpJLiqSG61MKF9TqfDVDJDbAJ1BqJFQ/tZ1U
4xaw+JekKw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZpIGfWiEBrG3Q+AWN1cRKeSOa/CDRdHr5NBYFH/IDhJ/Y1kjeN3kDbv/AbETrJnKGoU9EXN/2pUT
KF18zEDKoRrAeu/fv1ev6BfdXukihrRVgH3iSAu5c3WG5nTiEoAe8GgTHLguEMkU/gFk+RaGRnNe
AH+IWPK64N/cfhVZhhw=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bEbGnougkUJNEEp137e3KWyTp1SRyELmoiWnB1rmWN11lDaWBI/3Mk+Ax1nUdBNyIdVhcxj7m0B7
vUPGAb12ZYU5N4gxgAgD+tmnFl+SFvfR1JwPlrhqWMQ4wzGuALbjzkcXVht1tNLJ7d6gLn8IZ0zK
J1G826ATBadk3EdFXgU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Eg49/SbBigVS8KbFYYUAnUtZpnvmtXGBmqus5hcNYDVRIIiaRNtuR2Hbb3XbbhyKH0FZYs8pKARj
gAE7dz9GzM5E5ueMvO88tNOKOcqU4gF+uncWdlmHo3xl/COKMy0OwLFPp11NZfJB63PCWjAk1En3
+jy73/yAb53rwKHqNjE6AthGeUH0NdLFNdeBkNQx5EY2ugWegeL4iIIHM12owBtEdkojvTbJixbe
ilczKL50RkaSqWvN3gadF/O03BcufJSS9N80eJKHfIZ7Yqqj1rgbo3gB5wpY81niZC9eU5HWOpVs
u4XOqkSBIe+dgfxg0nNwhDfKTsH99LtnNRAx/w==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sDapw0WsH+J9ZoBenouuTES3qobkA+OlBh3ZC0TYJnYiF/o57VoTp0mj/jGyzpe4tDlc2H4HC6Fu
dcpxS2cNsKXipXnConEBfto+swfKSCYa7LnS/sYp6Szmd/KGrL9RwEsXjUmtAvlekEb3xUA7F73B
wh+TREr4452XHgEQOiBdHbc2/PA4qVkXtrExaXeZWtyAkCip0/0LLGEcuL4sWklgoIRWXOliTS9T
kOHl1r6lQjFOQhbNL2JBaf9rjo4CeJo9gMb3+20QclxYa5ek9v4olaPLGmuVdVshZcmkpia6wNsf
qpJ1dqLGIK1pMaBTuu5cLC/F8cGfxB+wE9jI3g==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uRRk4Q24ZeAWyuWLpEGFpeLvr739ht+7/2t3+kLJhpVwomZBbvl6K6a1+Lz2cAdAMs2TOzN3/fUA
i74LKe8jUulMgHJObWaljO29OoxtnKYPjK3S/rsQv3dEnOOKcol8QFz0cxYygoHR0ZhdSp1mBE2u
wX0CMZzZHoZelMuylsmPp2ZLSl2LVikF20g2mbMDO3YBt6mFxtrFgwrmPQ3nJxuyLjus/Nt/+OCe
R11QSgZbTzMyVkFV+MJOcbykbwugjgVwbNHbuukhf+Drz0KMgLmrL7m2Z0ZQW1NGh70dUhXCs87N
AX6MIxEk76/M1ZTkVqpDA4sGDOZBmmAE3a0gbQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5904)
`protect data_block
68hqkOrNlqcHe9GPJN1cThLONEzJKNGlcjdXYtvWQU2edjD3fk5XW6fIs2Fv7Er1pxJKQZFUFGDL
HKqOYuKU472t5I0Zh6ccW4is8lSXCjHHLLHV905XjC0vPI+nInsbrhPHsLTHVhqf0z6o+1Sa+/f9
3bOzo/AkKEqP/stG9xCVjmAVPY7tcF684i5Ao+pdp1j9To06r3V6Pkybj9D7VRuUuSazYGYK4KWK
g9WZN3AhkhQYI5guk/RhFfp7cxmrPth9DqbtMFkSvNoK2Yeo1IO4ULmQZAEGJTOMrvjRF39NriYB
ahw9Uqcq4KNG+6Q/+r0GLoXnVJPS9sPP0G4TOQnK7YTWYX0jxPhoyyy48d2E4Z92TVlby6BmMXTE
iCGskvkxxHh6+djpqz+QPMQjd1qsW8/o3pZzikxzDuboyGxoi29/EF3AB0D+UFsfj0rIHEPEKOeh
U3PqlJKIM+Hc/OmktnX6EtG8lGvVBrJn4+FcS7E+jteRttidsLiCi6pfyAJoheAivyFp1ZMkoe+9
Aj6XqzBwy/UEBtUFSlapyXDqzb2t1cU3AxQ0QhdqL3ojL5a9bvtuLk5GSQ5yyP6V473Unp97ZrWB
qU30dOgQ1dtfNxDO1jAU2vrO3IklFxWTokqE1xl1d/Sc+++7MhHNMOB+WOmH+sKfo0/a4ki83RYL
QfeBrhmrKBBsverFlbPBJLriFyqgvxyvaWObXtX+siSBuzL325HC8H+7g+kcL6PE+CyL+14yMhog
yT3GqrxAhw1/8j1X9SbUu7+VBWdz7gFvr/jvS4jwsWllSd1PGyeo0kzMvvhOfTe4RMj61kRsfd9d
ROPHoP8/f/zvVOcPo6zq1dCId4bs0wfM1oYGUTroYJAGDoHz/RhhNEim0CWK7WKsGoCoa0uIWk3Q
8k2bjADnsJ3tcSEtx+072smUcW8ZTZjZ3gSZ9605srkFFpLQFJIQX4Y8q+4AvIzTGOJPKdw6OC1v
8BiHQcho2DVX17mGQqWOMGpRqTmYDh/Uixk1FjhuGN1tvQLPAiN5wa/6eqA1vv3reA+NJhS2SfQ3
KFweQ8hoisKqnJ10aqD3bRTgkaliUqddZL7jRlZ74Bs6enyhzCMaNfvetIPLqVz25hsSCmI8njmq
MmgdwViOOavHMnN6tlnXok/6kC80I5juLikUqz9scyKvIkpTGKx59n+TjkKXn0CypsydrQmP+5b/
UcoEA0LvfENqj+I3j/VcV7+GgIQBAPQ/olVyIJlOUeidS7VMK9SWoRvFHc33duKiKQdkHLmGyRxs
sfvHJLuhFPjj9OF5fOuWXvi8YhIuFL470xIEh4JUW7JnKL9kkt6Ank2kUCERO1dM8H9caVf7EMWG
/Mc6vfNtF6PJ7RurOMCHEwmjHCRJjwJWyRFHLfIWeS7NvytvLiXfmS4Q3oh6N5T2WUIQfiCVdniD
nas/A5MeiRI/tHCoV6b554XWSDSAZ1mTW9QPLqI49AV1EKnCRtixqD42ir1PPcngSPayWPSZMypz
sRaGq0vDpv8RytSlChox+23Rb1EtGzt4mBI0/rIbywCmadFzeiiODqgEMEmdLIclL8kVb36OFXyY
ThdjPyUYk3ybVDLsCgQb6JLVaLB6vczUtCLtlCoSI56a+HD6ocYSTqaerSj+d3MvQqut1T+jkx5Z
GkmtydfGma5mI1VgdxB7o2dxYvx8xDuDTuDBDcVu9Z7V+O/Rfav1yv2XM/mYJTzXehbuxAXxoUI4
1/dGfjTmHves0KUAdFIspXqs7QVqn8HrQhm1quGFKcyjQ1DpQ8ZhvibLczcPFM5ISbqtctpM5fYZ
CDPZhV9dVRoD17usqXRZoBMC8GsGziqzBlxEC4NOXjrt5YupozxGnCMXh9PngpsiSW3dustU1HFj
A5hxUG/7L1u8SZoXSacqqMy0z98PaMPo5x27g12MRzR2sMUxXVNeORfVAWFRrmiEjKDkTWwWkoKz
vohzNWVR4oIF8o5+31SNTCoPTB0yuvVVEQpBZMH3xv6Y/1oFxq1OnBpOrcT0gNH/goS/cxwHvNaS
OXfOzf5KtM20MOEFyFZt+2sKrd/VQeMRYV90DQmx0l3F6cILV7GReGaTAHJLx9Zl+lv8gk8aF3g9
98Z9H0apb8PjaPeBM9vCQVYDYUppPOlqOGAFVW/KnQ3eKiQ+oDOOf1iretV+CtFMsDCFDGIo3asL
yHkMVaTxBLImBQozbaJd/3WaBXr3tgsTNuLokWE5NG+postfcuGdcaBBRx+CFtmR+6MgE+7NaLZ4
00ZNm8n5tkMX6vWc1bDy77m+hNohMFp3Sf3qyJthXfCPQHzbCG0RUr1VhkWZgw18iDaZeAkV+aGJ
X57VfKZ3sjVwqqByZeULYjJB+o4x5Zx+EjQ23Q5uLd9ljbnCKGZ5LzGS0UXmSnhwwZXYZiR7pKii
W1FDmTUOpKf0o5yPmy80PMyaF4eaq0USjzv/1cgitCu+f53zRGkcJYnNqYFXtOKRPnB28mv076g4
dj+r4H/L0EJwfeeg4hVu6kcZNYPjJjQVMlsSHS/FCp8wUsLIFubetlL4JOMP3W3fm/0Ku1d+IG7a
B8o2lWifLNo5J6MY3N2J6nZGK1PYsJKrLayVwflXDQ+cY1JpY8sVbmbwu0g0NvRFN16lktap4/cp
xNpoPAFkIS4PLJTaqBpbP/Wcu4344Bmnd5fWLj3J98qQL4wKqzh6/mwzuDG/aZ53m/9YmZLK7g6/
Z3IgQBaTJEeM7mB8tuDxulXzK6sq23M44NlVVEGhbKraDQBZZha37dqigs4i17hSUJm91hyziprS
US58qYrBWty5WpvhODnrqVrcohaqdaltlTgKcjz+wcc3vbYOKXevBwkIH0zA3/TaNKhrbab7zcc1
Hum8aSldMIStLclSIBzWIyyRL12cOCqbdu4Frcn6wHMrCUe+1R+fJTtPeAokxXAQ3lVv/yYPoo3I
8Kh8bd/PBJPIA2vAl1QNSUasnsBhVzRqLrZsE9fmcAQoDN05SqCtuD+1qurvR0ljuZoGJO+EhI+o
vBmtgxJTx7SFrFMCd6j3/VWog8bQoUnMCh+m2aRiP9JfsU/KfaxdmwAiJtKZjCdRCHFHsmnwBbuR
JjnnnDfa13pmWoHAiRxptj5vzud+vvBUUIUi+b9ZW/YX1yF+G/12JTgQI4PhyhifKyjwTT/8TjcJ
zJgxNCClVs2kVi9bRyVPFjIajw4kQkn+sl6+xDprLFbf9PLwPYit5uP9CKkE/rT5UujxFGSonMU1
UVEGXhWztFloKMnptBYSiAGDL7UmA4HLCEFTynbg9zg0yEOrcnEgJyshieH9zmDl1MfOtckBhMhS
pXaSFJEadPDg4bMJ2MSNSY/1+ndgNQ0zyP647YzGX5ZXrl1NeoOmgKpN/iKQVV69sUkjycQ+EbQh
hquqGpnINm5qd4AWjS5PS6qFi+oeC312ZCZlt1OYho2ZwsbxXHN4LRpbxABnBsiCuyeoYYNPwE9Y
kDdse526cUZMUjTu+jUmYIkja7N/CvM3ExNe0Ij589f6rmW1u65yU2WZEeW4BqfC5qidD1Gx/4ji
w0N3inTXJnHaDXK0hoQAmGO/cHdr0HVj09tZkUodJ9AOjFizbt0pRFgirYxo2cWoxnlc28NtoabI
fM6HfqX/xEQXPiYhWI5TtZ6hZ5y7iN0s9dwBqPsJfMq2VE4EAPQubJ7VNzwLQsnjwzPNuyo3JqN6
vNni2NaYwXbwoA0yhVq8DS0i25bAGHr79mF5BTv4RFKfEsz1e8IJ7Ogm5Ln3L8/J01xyqjcZ3auo
EygjfG+tCPMAP2UsITGZE7p/QIaYgMyING3ozLkfCErCeaZ5toY7ghpAeYKZCQ+1gWF+NJVgVVew
M5Uftn6s+UfhO3WsJ2d+Y6zZBry7AMJT3BnaX5lkvcXNbc1v0TbdXbnLFnc0BsClUKEBDM0ifdq4
KpLOhvEU98WOVFEOW0F9VlMBRaPv11i5OjMPeTCbFqNKtKrCuckjOD1gl1AK6pHr+rRugLf1p6mS
PeWj2dtREwF0GBoJO1n+2ruwtS+zJwAxYL5BRb775Y9QIZta3BW5zgXmO9vq+5YBtht4RNS5ZhHk
D6htw2HnASrXVW6vtYMq9YsiE3Hyx/EPLAR4u09Ncq/lGIZ88M3YjiEthQGv4U2bIxZFTHAc/+Qi
Emu4/mYju4MvlBTRBlBBNk4YFm9X9P8IhgII6dw35qERH0H81dxDC4EgXEIukwKisQ3WZUeXGkeG
gRzhsiEbtQDn9L4bvKjzQYWZWGGq5McbxjbiHaBErGgj7NWlAYfg3hvSHuwVHCw4JJ0xH0dxF8KU
ymz+8JE9PQmPfrcM2Yy37vY2ZuQcY2e/SH+ccbQ7J2TvKE/kMqpw5NCpcFVK1B9LhbzGnIzEkb6f
3+t7ZK6lEvbRmgjr8HTxSBUi7AD9+t56O0E+48raWfKmrk58v7rkOcmZ9b8IhJGcibNDZhcbWB4w
QNnW0UZ8JiAt4tyEVu+ZpTb9u6p6zxmuZv6tryUw47/yhB4q/RTPO3WoXLL2A8EEgFDkPw37Gccp
CkPyGHDVxKbVwYvbnOlKRLVSMpZZ5LVwhGZQPgIpbNbMKy05eplOoxJHv/1lktIzGmaM9Kwh769V
n2EDalNn34WbD6M2qVQ4sc2l+Y2kkMk/c+6TuJGp/G+kRMiwzlJgVIUPUtzgYswjfSVxJgyeOO0R
K3deDCbArgZigKobgTRCzopqZAd6OAmZ4fGPzI7tGFq5hky5TMVv8Xlfn/RbM3Nf092PPKLGqyZu
BDmqkmcYCKOYsLT793n99SG3CC9o7nIL/CghuSx7BlEN0cllzuXlMLoa1Up1qBWhF0kj3bmfMlDx
IoKqhu/TQ+JHD7yxsFPoiJ6AMsaXkecXbgd6vW5KQ90QmP1UcyEiROMHOA6Yjkc5oqAy434gXBx6
sjF0Lev2Gd+RvRnIiTltCwWavxd/v6YNe9NY8htmMBZQfhYNp3fre/bkY/WzuZ5Kdp6s4QRdrir/
LEY5ZvJDn2UPr2wkKtgRds+aIgWouEYvHL3PbwEQXSQwQpEcoUF79EIV5KL/8lshQnVuGHFgVJ7U
diCCIk4+RngiuTN1XBVI+NRCalhYydD50yV33J+VVNa5WFhVHxJ4Fbjz89n5mRBtvVbypqQlyAqZ
RS52HMMrysP4fWIOMlH7E7zjezb8sMGUXO3nPy02wJxnbXYimHblxfM60FSa1GuZhC6INGnzZptI
2usg0hBIppIzuGBZ434xC97YpoLVs3fydKkgf7UyZWHpi75x8Ol7SFxRnLGUnJ48i4GP6pyiZLBt
PoR7sMrRXqVRDPOG39a3V0B281YLmlmSA8FK25NAlvtsNlC/0Neg3W6GjiCLFDHsCo8IwNAZUdcu
QcHMsP03N8xwIJh9+BkhCXO6XrC5d96d6MoNx9d9IoP0sKrSC8bZzRgGd330am7jF0IMsEjNae2U
AnQSAHH3WD0MWr3dFy+/VhEVbrl9/3b+EJQm92ViAn9pJGxEStZrrVOWf81BdLhUkATId87+302W
1B31ZNjeQBeFHhsZA2ziSO/HsgAItaD0jpayrC2AgRJ0yA2u5HQcQJR1mYOYQSbxl30mv4Diu3Z+
a/xxh3Bphuarz+cY5mKMeg2KgjfTfn2O5nEPTIcMFsLpHApTm1Jh4eVvaGVXvUYY8By5ulbZ1o3X
1pk/VJzGJnVTST7N7wWDCuYuBOeIDuCiBoCbtVosPzICLGVpJY29jZdlP7Y40yBfIrWpIMZ9G1NT
Nnxi19JomECba3GxjQfncgfNxTeXyx29KkIqWlnct2kZp8k+R3jgRmllMRlaZ/xsL5ioEMT+ekcV
DWu7Nh6kQ8gP8F+NLj8VjReZmJBz9kMwmWrtR1kEMIpmYI1Y5CpBbp4wEBiW6KmeQnbcdOg0750H
f4jc4pe5k1ABuTOER2FsV97S1HedabQtlYFdgSZxCchCt/sjOJqd/QjwghPxni0oojvZUhCsHH3i
6ASov4Nv/M9WFWeI5t86dOTg9IVOv9usqSqfUwbsEpOyG0cBAaO13Nt8UchPEXAn1C36HSfNu/Ua
h7DqsB8XhNCaiXWFfcYsySM3Jh1xVVEZUznaL7djQiQs5N8mS5zOL3kPjRjZ+oDMAyuE1GR65g7u
LbSvFR9RzF2bI06WaAVH20diV5Y/aYNOcuxtV/2essVNv6Kdu0XjWzUbXIGx6GzcYB1HjpKTuwo3
mMEjQI8ZN8+QBy0L0oIzbX4H9ZVlk6xzbidOHhAyIX3F03J82qTiGiFoGwi5cy3FGi8dFjfnl1gi
2icO/8+xOpPU3odQeaEBWCH5aVD9rLvrYTbs2xJPCNaU88PRrbiaicV1xYAkX7TjRGH6rrYdLypR
aG45W7tpHgzDLiDKePxwXU97O0e4Szma/qzCYT3BZvCNo6RmxdIxnhkgMkcCb1b8xkaccGZxOw8T
056BF+I1qLD/Qrb9+rCD1dS3oymdgZN0jALHJUD1bbJve1BEG2XdPof/ZyeqS/VM3GAyuJ7puU+f
t217cY0nTJLH3b6FEdcZdoxVIKHqTLNkqmwvURjcMGzPI3r1I3plBrQrtBs5EzjhT3fyW3tkwsur
CaWLd5zazLmETZTUsy5L2x1g7tkl0usMNo368CqjOFtOPh2yJ/s/V/6bG3FdiC9L0qk7TGA/+wbl
pYhig639pwuqogDE2FKWsg0t0afrDc9HnPMS6isSCryEb92r89tzcJ3dfjTPH+fJTCropM5rQJ7o
KCPDLb9haeWQfNp9xRAFKuIZ3Q15is69qC/G/Ni6TnmyjdmTmQ8YQPWE5nZH7Yt+dmt+cImbwxIQ
3VS4uCfNY8JhCRbUs/i6iVhBxvXVwIsIKYQkKtoRRyil4dAmj97fsvrdTR2s8Uu3zohrWGwuz4Ef
ljYnMYCfoOzXKvvPzsEFrkR+XH5PulpuHAyBwT104jcon5l2WB2F2JaEcSRuu+QHXw6N22FQ06FQ
N16Ms0KPFdpQD5zMRtD5IiMGWP19FJnJ1QRw/AJsu09z63Kn/BXVCwXH9gkIINl5E8LBK1oF8Fha
n2UkhF4jZdTNEKoMgV9pus5P3cB/pcXx5bj4i5m3ocJRM1X6ZdEwcjSJww88jADc5UhTIH8ZP+/S
cY1CMG4F3GXsihsb7E1lwK1BXeNRCKZn07kWDQD0w5zfk4B0b4o9Re5TB2DWfUAlPCFQoZuEIV/5
QuYNgj/h2+M6kSOuXAwiR9PVZDgnKXOo4BU1/jg1E0na9qe9r9WNtVAOx40H1Oz8EKTc9ygp/9rZ
hm5khAfCeZ2jIKk9XDK2b7ZAG0qAsGLduqIiULS6spFU+3JochhYiG5s6sCnxUNkGjgsmWMG+OqX
WlAfoIbfAdESgw9ooS84iyieBGXdB+Ff3GcweVtVfhHW9ARkDGws6LQdYSwLUNsMm2yztf3U+D6z
+Dt+eyKcwPl4Jp22aoIboo11408yqTf65yd+6rkCUZNvNCyjJv96Yc5YbpaTOmNp37tFm8HFHBiT
jUgoRLZ3623nuoNN6hDiIftcyGHvyvcfSauYfZ9qXy6+bvm/AWK2uFsoMvzWKzYS4MkienQfxTwH
lgze0FkqwIjb7iaMuRiSFY5ZNiPGiiKwFrn96mzjWWcWySIQfz6DrHy2V1rhaUgbJZaNx6Xz1RWT
ALp49eaki33RXxI2u022xQ0qPfqizXqsbN1l8Qi14ch2IlqsHMOCrcl+VH9ese+SNNLyN1kQCGpU
/y5WFHpm4p4qFM+5z3lsSPyjW7CaFrurIjpbYx6qT7abRYi2NHW6G5IbbUIzqhLJB4FzAezPnnRe
h4yl48wgFNYGRBNOZEI4+3nnjTO0+cTFheq+8fkTqLJW
`protect end_protected
